
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_aes_dec_KEY_SIZE2 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_aes_dec_KEY_SIZE2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_aes_dec_KEY_SIZE2.all;

entity key_expansion is

   port( KEY_I : in std_logic_vector (7 downto 0);  VALID_KEY_I, CLK_I, RESET_I
         , CE_I : in std_logic;  DONE_O : out std_logic;  GET_KEY_I : in 
         std_logic;  KEY_NUMB_I : in std_logic_vector (5 downto 0);  KEY_EXP_O 
         : out std_logic_vector (31 downto 0));

end key_expansion;

architecture SYN_Behavioral of key_expansion is

   component IVI
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component EO
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NR2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EN
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component ND2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AN3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component AO7
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component AO4
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component AO6
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component AO2
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component EOI
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component ND3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component NR3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component AO3
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component EON1
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component EO1
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component NR4
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component IVDA
      port( A : in std_logic;  Y, Z : out std_logic);
   end component;
   
   component ND2I
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component ND4
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component ENI
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NR2I
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AN2I
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AO1P
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component AN4
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FD1
      port( D, CP : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal v_KEY32_IN_31_port, v_KEY32_IN_30_port, v_KEY32_IN_29_port, 
      v_KEY32_IN_28_port, v_KEY32_IN_27_port, v_KEY32_IN_26_port, 
      v_KEY32_IN_25_port, v_KEY32_IN_24_port, v_KEY32_IN_23_port, 
      v_KEY32_IN_22_port, v_KEY32_IN_21_port, v_KEY32_IN_20_port, 
      v_KEY32_IN_19_port, v_KEY32_IN_18_port, v_KEY32_IN_17_port, 
      v_KEY32_IN_16_port, v_KEY32_IN_15_port, v_KEY32_IN_14_port, 
      v_KEY32_IN_13_port, v_KEY32_IN_12_port, v_KEY32_IN_11_port, 
      v_KEY32_IN_10_port, v_KEY32_IN_9_port, v_KEY32_IN_8_port, 
      v_KEY32_IN_7_port, v_KEY32_IN_6_port, v_KEY32_IN_5_port, 
      v_KEY32_IN_4_port, v_KEY32_IN_3_port, v_KEY32_IN_2_port, 
      v_KEY32_IN_1_port, v_KEY32_IN_0_port, v_CALCULATION_CNTR_7_port, 
      v_CALCULATION_CNTR_6_port, v_CALCULATION_CNTR_5_port, 
      v_CALCULATION_CNTR_4_port, v_CALCULATION_CNTR_3_port, 
      v_CALCULATION_CNTR_2_port, v_CALCULATION_CNTR_1_port, 
      v_CALCULATION_CNTR_0_port, i_SRAM_ADDR_WR0, i_SRAM_ADDR_WR01, 
      i_SRAM_ADDR_WR02, i_SRAM_ADDR_WR03, i_SRAM_ADDR_WR04, i_SRAM_ADDR_WR05, 
      v_KEY_COL_OUT0_31_port, v_KEY_COL_OUT0_30_port, v_KEY_COL_OUT0_29_port, 
      v_KEY_COL_OUT0_28_port, v_KEY_COL_OUT0_27_port, v_KEY_COL_OUT0_26_port, 
      v_KEY_COL_OUT0_25_port, v_KEY_COL_OUT0_24_port, v_KEY_COL_OUT0_23_port, 
      v_KEY_COL_OUT0_22_port, v_KEY_COL_OUT0_21_port, v_KEY_COL_OUT0_20_port, 
      v_KEY_COL_OUT0_19_port, v_KEY_COL_OUT0_18_port, v_KEY_COL_OUT0_17_port, 
      v_KEY_COL_OUT0_16_port, v_KEY_COL_OUT0_15_port, v_KEY_COL_OUT0_14_port, 
      v_KEY_COL_OUT0_13_port, v_KEY_COL_OUT0_12_port, v_KEY_COL_OUT0_11_port, 
      v_KEY_COL_OUT0_10_port, v_KEY_COL_OUT0_9_port, v_KEY_COL_OUT0_8_port, 
      v_KEY_COL_OUT0_7_port, v_KEY_COL_OUT0_6_port, v_KEY_COL_OUT0_5_port, 
      v_KEY_COL_OUT0_4_port, v_KEY_COL_OUT0_3_port, v_KEY_COL_OUT0_2_port, 
      v_KEY_COL_OUT0_1_port, v_KEY_COL_OUT0_0_port, i_INTERN_ADDR_RD0, 
      i_INTERN_ADDR_RD01, i_INTERN_ADDR_RD02, i_INTERN_ADDR_RD03, 
      i_INTERN_ADDR_RD04, i_INTERN_ADDR_RD05, v_TEMP_VECTOR_31_port, 
      v_TEMP_VECTOR_30_port, v_TEMP_VECTOR_29_port, v_TEMP_VECTOR_28_port, 
      v_TEMP_VECTOR_27_port, v_TEMP_VECTOR_26_port, v_TEMP_VECTOR_25_port, 
      v_TEMP_VECTOR_24_port, v_TEMP_VECTOR_23_port, v_TEMP_VECTOR_22_port, 
      v_TEMP_VECTOR_21_port, v_TEMP_VECTOR_20_port, v_TEMP_VECTOR_19_port, 
      v_TEMP_VECTOR_18_port, v_TEMP_VECTOR_17_port, v_TEMP_VECTOR_16_port, 
      v_TEMP_VECTOR_15_port, v_TEMP_VECTOR_14_port, v_TEMP_VECTOR_13_port, 
      v_TEMP_VECTOR_12_port, v_TEMP_VECTOR_11_port, v_TEMP_VECTOR_10_port, 
      v_TEMP_VECTOR_9_port, v_TEMP_VECTOR_8_port, v_TEMP_VECTOR_7_port, 
      v_TEMP_VECTOR_6_port, v_TEMP_VECTOR_5_port, v_TEMP_VECTOR_4_port, 
      v_TEMP_VECTOR_3_port, v_TEMP_VECTOR_2_port, v_TEMP_VECTOR_1_port, 
      v_TEMP_VECTOR_0_port, N1748, N1749, N1750, N1751, N1752, N1753, N1754, 
      n13, n15, n16, n17, n18, n19, n20, n21, n24, n25, n26, n27, n29, n30, n31
      , n32, n34, n35, n36, n37, n39, n40, n41, n42, n44, n45, n46, n47, n49, 
      n50, n51, n52, n54, n55, n56, n57, n60, n61, n62, n63, n64, n65, n66, n67
      , n68, n70, n73, n74, n75, n76, n77, n78, n79, n80, n82, n83, n84, n85, 
      n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, 
      n100, n101, n102, n103, n104, n105, n106, n107, n108, n110, n111, n112, 
      n113, n114, n115, n116, n117, n118, n119, n120, n121, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n164, n165, n166, n167, n168, n169, n171, n172, n173, n174, n175, n176, 
      n177, n178, n179, n181, n182, n183, n184, n185, n186, n187, n188, n189, 
      n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n201, n202, 
      n203, n204, n205, n206, n207, n208, n210, n211, n212, n213, n214, n215, 
      n216, n218, n219, n220, n221, n222, n223, n225, n226, n230, n231, n233, 
      n239, n240, n242, n243, n244, n247, n252, n254, n256, n262, n263, n264, 
      n266, n267, n268, n271, n273, n274, n275, n277, n278, n279, n280, n281, 
      n282, n283, n285, n287, n288, n289, n290, n291, n292, n294, n295, n296, 
      n297, n298, n299, n300, n302, n304, n305, n306, n307, n308, n309, n310, 
      n311, n312, n313, n315, n316, n317, n318, n319, n320, n321, n322, n323, 
      n324, n326, n327, n328, n329, n330, n331, n332, n333, n334, n336, n337, 
      n338, n339, n340, n341, n342, n343, n344, n345, n346, n355, n356, n357, 
      n358, n367, n368, n369, n370, n379, n380, n381, n382, n391, n392, n393, 
      n394, n395, n396, n397, n398, n407, n408, n409, n410, n419, n420, n421, 
      n422, n431, n432, n433, n434, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, 
      n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, 
      n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, 
      n524, n525, n526, n527, n528, n529, n530, n532, n533, n534, n535, n536, 
      n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, 
      n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, 
      n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, 
      n573, n574, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, 
      n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, 
      n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, 
      n610, n611, n612, n613, n614, n615, n616, n617, n618, n620, n621, n622, 
      n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, 
      n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, 
      n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, 
      n659, n660, n661, n662, n664, n665, n666, n667, n668, n669, n670, n671, 
      n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, 
      n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, 
      n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n708, 
      n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, 
      n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, 
      n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, 
      n745, n746, n747, n748, n749, n750, n752, n753, n754, n755, n756, n757, 
      n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, 
      n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, 
      n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, 
      n794, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, 
      n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, 
      n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, 
      n831, n832, n833, n834, n835, n836, n837, n838, n840, n841, n842, n843, 
      n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, 
      n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, 
      n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, 
      n880, n881, n882, n884, n885, n886, n887, n888, n889, n890, n891, n892, 
      n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, 
      n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, 
      n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n928, n929, 
      n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, 
      n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, 
      n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, 
      n966, n967, n968, n969, n970, n972, n973, n974, n975, n976, n977, n978, 
      n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, 
      n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002
      , n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, 
      n1013, n1014, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, 
      n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, 
      n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, 
      n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, 
      n1054, n1055, n1056, n1057, n1058, n1060, n1061, n1062, n1063, n1064, 
      n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, 
      n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, 
      n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, 
      n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1104, n1105, 
      n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, 
      n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, 
      n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, 
      n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, 
      n1146, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, 
      n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, 
      n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, 
      n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, 
      n1187, n1188, n1189, n1190, n1192, n1193, n1194, n1195, n1196, n1197, 
      n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, 
      n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, 
      n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, 
      n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1236, n1237, n1238, 
      n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, 
      n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, 
      n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, 
      n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, 
      n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, 
      n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, 
      n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, 
      n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, 
      n1320, n1321, n1322, n1324, n1325, n1326, n1327, n1328, n1329, n1330, 
      n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, 
      n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, 
      n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, 
      n1361, n1362, n1363, n1364, n1365, n1366, n1368, n1369, n1370, n1371, 
      n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, 
      n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, 
      n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, 
      n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1412, 
      n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, 
      n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, 
      n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, 
      n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, 
      n1453, n1454, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, 
      n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, 
      n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, 
      n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, 
      n1494, n1495, n1496, n1497, n1498, n1500, n1501, n1502, n1503, n1504, 
      n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, 
      n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, 
      n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, 
      n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1544, n1545, 
      n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, 
      n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, 
      n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, 
      n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, 
      n1586, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, 
      n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, 
      n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, 
      n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, 
      n1627, n1628, n1629, n1630, n1632, n1633, n1634, n1635, n1636, n1637, 
      n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, 
      n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, 
      n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, 
      n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1676, n1677, n1678, 
      n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, 
      n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, 
      n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, 
      n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, 
      n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, 
      n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, 
      n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748_port, 
      n1749_port, n1750_port, n1751_port, n1752_port, n1753_port, n1754_port, 
      n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1764, n1765, 
      n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, 
      n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, 
      n1786, n1787, n1788, n1789, n1790, n1791, n1794, n1795, n1796, n1797, 
      n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, 
      n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, 
      n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, 
      n1828, n1829, n1830, n1831, n1834, n1835, n1836, n1837, n1838, n1839, 
      n1840, n1841, n1842, n1845, n1846, n1848, n1849, n1850, n1851, n1852, 
      n1853, n1854, n1855, n1856, n1857, n1860, n1863, n1864, n1869, n1870, 
      n1871, n1873, n1874, n1879, n1880, n1881, n1884, n1885, n1886, n1887, 
      n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, 
      n1902, n1907, n1909, n1911, n1912, n1913, n1914, n1915, n1916, n1918, 
      n1919, n1920, n1923, n1924, n1925, n1926, n1927, n1928, n1930, n1932, 
      n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1942, n1943, 
      n1944, n1945, n1946, n1948, n1950, n1951, n1952, n1953, n1954, n1955, 
      n1957, n1958, n1959, n1960, n1961, n1963, n1964, n1965, n1969, n1970, 
      n1971, n1972, n1973, n1975, n1976, n1977, n1978, n1979, n1980, n1983, 
      n1985, n1986, n1987, n1988, n1990, n1991, n1992, n1993, n1994, n1995, 
      n1996, n1997, n1998, n2000, n2002, n2003, n2004, n2005, n2006, n2007, 
      n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, 
      n2018, n2019, n2020, n2021, n2022, n2024, n2025, n2026, n2027, n2028, 
      n2029, n2030, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, 
      n2040, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2051, 
      n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, 
      n2062, n2063, n2064, n2065, n2067, n2068, n2069, n2070, n2071, n2072, 
      n2073, n2074, n2075, n2077, n2078, n2079, n2080, n2081, n2082, n2083, 
      n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2092, n2093, n2094, 
      n2095, n2096, n2097, n2099, n2100, n2102, n2104, n2105, n2106, n2107, 
      n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, 
      n2118, n2119, n2120, n2122, n2123, n2124, n2125, n2126, n2128, n2129, 
      n2130, n2131, n2132, n2133, n2135, n2136, n2137, n2138, n2139, n2140, 
      n2141, n2142, n2143, n2144, n2145, n2147, n2148, n2149, n2151, n2152, 
      n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2162, n2163, 
      n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, 
      n2174, n2176, n2178, n2179, n2180, n2182, n2184, n2185, n2186, n2187, 
      n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, 
      n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2206, n2207, n2208, 
      n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2218, n2219, 
      n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, 
      n2231, n2232, n2234, n2235, n2236, n2237, n2238, n2239, n2241, n2242, 
      n2243, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, 
      n2254, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, 
      n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2275, 
      n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, 
      n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, 
      n2296, n2298, n2299, n2300, n2301, n2302, n2303, n2306, n2307, n2309, 
      n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, 
      n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, 
      n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, 
      n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, 
      n2480, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, 
      n2493, n2495, n2496, n2497, n2498, n2499, n2500, n2502, n2503, n2505, 
      n2506, n2507, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, 
      n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, 
      n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, 
      n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, 
      n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, 
      n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, 
      n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, 
      n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, 
      n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, 
      n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, 
      n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, 
      n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, 
      n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, 
      n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, 
      n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, 
      n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, 
      n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, 
      n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, 
      n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, 
      n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, 
      n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, 
      n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, 
      n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, 
      n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, 
      n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, 
      n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, 
      n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, 
      n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, 
      n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, 
      n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, 
      n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, 
      n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, 
      n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, 
      n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, 
      n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, 
      n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, 
      n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, 
      n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, 
      n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, 
      n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, 
      n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, 
      n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, 
      n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, 
      n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, 
      n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, 
      n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, 
      n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, 
      n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, 
      n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, 
      n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, 
      n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, 
      n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, 
      n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, 
      n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, 
      n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, 
      n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, 
      n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, 
      n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, 
      n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, 
      n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, 
      n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, 
      n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, 
      n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, 
      n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, 
      n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, 
      n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, 
      n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, 
      n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, 
      n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, 
      n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, 
      n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, 
      n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, 
      n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, 
      n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, 
      n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, 
      n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, 
      n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, 
      n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, 
      n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, 
      n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, 
      n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, 
      n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, 
      n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, 
      n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, 
      n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, 
      n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, 
      n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, 
      n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, 
      n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, 
      n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, 
      n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, 
      n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, 
      n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, 
      n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, 
      n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, 
      n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, 
      n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, 
      n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, 
      n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, 
      n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, 
      n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, 
      n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, 
      n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, 
      n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, 
      n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, 
      n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, 
      n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, 
      n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, 
      n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, 
      n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, 
      n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, 
      n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, 
      n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, 
      n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, 
      n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, 
      n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, 
      n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, 
      n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, 
      n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, 
      n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, 
      n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, 
      n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, 
      n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, 
      n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, 
      n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, 
      n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, 
      n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, 
      n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, 
      n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, 
      n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, 
      n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, 
      n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, 
      n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, 
      n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, 
      n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, 
      n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, 
      n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, 
      n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, 
      n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, 
      n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, 
      n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, 
      n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, 
      n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, 
      n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, 
      n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, 
      n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, 
      n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, 
      n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, 
      n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, 
      n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, 
      n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, 
      n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, 
      n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, 
      n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, 
      n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, 
      n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, 
      n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, 
      n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, 
      n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, 
      n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, 
      n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, 
      n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, 
      n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, 
      n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, 
      n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, 
      n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, 
      n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, 
      n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, 
      n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, 
      n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, 
      n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, 
      n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, 
      n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, 
      n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, 
      n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, 
      n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, 
      n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, 
      n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, 
      n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, 
      n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, 
      n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, 
      n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, 
      n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, 
      n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, 
      n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, 
      n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, 
      n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, 
      n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, 
      n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, 
      n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, 
      n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, 
      n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, 
      n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, 
      n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, 
      n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, 
      n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, 
      n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, 
      n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, 
      n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, 
      n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, 
      n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, 
      n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, 
      n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, 
      n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, 
      n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, 
      n4557, n4561, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, 
      n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, 
      n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, 
      n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, 
      n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, 
      n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, 
      n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, 
      n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, 
      n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, 
      n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, 
      n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, 
      n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, 
      n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, 
      n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, 
      n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, 
      n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, 
      n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, 
      n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, 
      n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, 
      n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, 
      n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, 
      n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, 
      n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, 
      n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, 
      n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, 
      n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, 
      n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, 
      n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, 
      n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, 
      n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, 
      n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, 
      n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, 
      n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, 
      n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, 
      n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, 
      n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, 
      n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, 
      n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, 
      n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, 
      n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, 
      n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, 
      n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, 
      n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, 
      n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, 
      n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, 
      n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, 
      n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, 
      n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, 
      n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, 
      n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, 
      n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, 
      n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, 
      n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, 
      n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, 
      n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, 
      n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, 
      n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, 
      n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, 
      n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, 
      n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, 
      n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, 
      n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, 
      n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, 
      n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, 
      n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, 
      n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, 
      n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, 
      n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, 
      n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, 
      n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, 
      n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, 
      n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, 
      n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, 
      n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, 
      n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, 
      n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, 
      n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, 
      n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, 
      n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, 
      n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, 
      n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, 
      n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, 
      n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, 
      n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, 
      n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, 
      n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, 
      n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, 
      n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, 
      n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, 
      n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, 
      n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, 
      n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, 
      n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, 
      n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, 
      n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, 
      n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, 
      n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, 
      n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, 
      n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, 
      n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, 
      n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, 
      n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, 
      n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, 
      n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, 
      n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, 
      n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, 
      n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, 
      n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, 
      n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, 
      n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, 
      n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, 
      n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, 
      n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, 
      n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, 
      n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, 
      n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, 
      n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, 
      n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, 
      n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, 
      n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, 
      n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, 
      n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, 
      n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, 
      n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, 
      n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, 
      n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, 
      n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, 
      n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, 
      n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, 
      n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, 
      n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, 
      n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, 
      n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, 
      n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, 
      n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, 
      n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, 
      n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, 
      n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, 
      n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, 
      n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, 
      n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, 
      n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, 
      n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, 
      n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, 
      n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, 
      n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, 
      n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, 
      n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, 
      n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, 
      n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, 
      n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, 
      n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, 
      n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, 
      n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, 
      n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, 
      n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, 
      n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, 
      n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, 
      n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, 
      n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, 
      n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, 
      n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, 
      n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, 
      n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, 
      n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, 
      n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, 
      n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, 
      n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, 
      n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, 
      n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, 
      n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, 
      n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, 
      n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, 
      n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, 
      n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, 
      n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, 
      n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, 
      n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, 
      n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, 
      n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, 
      n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, 
      n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, 
      n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, 
      n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, 
      n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, 
      n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, 
      n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, 
      n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, 
      n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, 
      n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, 
      n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, 
      n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, 
      n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, 
      n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, 
      n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, 
      n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, 
      n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, 
      n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, 
      n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, 
      n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, 
      n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, 
      n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, 
      n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, 
      n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, 
      n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, 
      n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, 
      n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, 
      n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, 
      n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, 
      n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, 
      n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6673, 
      n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, 
      n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, 
      n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, 
      n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, 
      n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, 
      n6724, n6725, n6726, n6727, n6728, n6729, n6762, n6763, n1, n2, n3, n4, 
      n5, n6, n7, n8, n9, n10, n11, n12, n14, n22, n23, n28, n33, n38, n43, n48
      , n53, n58, n59, n69, n71, n72, n81, n109, n122, n150, n163, n170, n180, 
      n200, n209, n217, n224, n227, n228, n229, n232, n234, n235, n236, n237, 
      n238, n241, n245, n246, n248, n249, n250, n251, n253, n255, n257, n258, 
      n259, n260, n261, n265, n269, n270, n272, n276, n284, n286, n293, n301, 
      n303, n314, n325, n335, n347, n348, n349, n350, n351, n352, n353, n354, 
      n359, n360, n361, n362, n363, n364, n365, n366, n371, n372, n373, n374, 
      n375, n376, n377, n378, n383, n384, n385, n386, n387, n388, n389, n390, 
      n399, n400, n401, n402, n403, n404, n405, n406, n411, n412, n413, n414, 
      n415, n416, n417, n418, n423, n424, n425, n426, n427, n428, n429, n430, 
      n435, n436, n437, n438, n439, n440, n441, n442, n443, n487, n531, n575, 
      n619, n663, n707, n751, n795, n839, n883, n927, n971, n1015, n1059, n1103
      , n1147, n1191, n1235, n1279, n1323, n1367, n1411, n1455, n1499, n1543, 
      n1587, n1631, n1675, n1719, n1763, n1792, n1793, n1832, n1833, n1843, 
      n1844, n1847, n1858, n1859, n1861, n1862, n1865, n1866, n1867, n1868, 
      n1872, n1875, n1876, n1877, n1878, n1882, n1883, n1888, n1889, n1890, 
      n1901, n1903, n1904, n1905, n1906, n1908, n1910, n1917, n1921, n1922, 
      n1929, n1931, n1941, n1947, n1949, n1956, n1962, n1966, n1967, n1968, 
      n1974, n1981, n1982, n1984, n1989, n1999, n2001, n2023, n2031, n2041, 
      n2050, n2066, n2076, n2091, n2098, n2101, n2103, n2121, n2127, n2134, 
      n2146, n2150, n2161, n2175, n2177, n2181, n2183, n2205, n2217, n2220, 
      n2233, n2240, n2244, n2255, n2274, n2297, n2304, n2305, n2308, n2310, 
      n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, 
      n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, 
      n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, 
      n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, 
      n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, 
      n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, 
      n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, 
      n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, 
      n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, 
      n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, 
      n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, 
      n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, 
      n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2479, n2481, 
      n2491, n2492, n2494, n2501, n2504, n2508, n4558, n4559, n4560, n4562, 
      n6670, n6671, n6672, n6730, n6731, n6732, n6733, n6734, n6735, n6736, 
      n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, 
      n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, 
      n6757, n6758, n6759, n6760, n6761, n6764, n6765, n6766, n6767, n6768, 
      n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, 
      n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, 
      n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, 
      n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n_1000, 
      n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, 
      n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, 
      n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, 
      n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, 
      n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, 
      n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, 
      n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, 
      n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, 
      n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, 
      n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, 
      n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, 
      n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, 
      n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, 
      n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, 
      n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, 
      n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, 
      n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, 
      n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, 
      n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, 
      n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, 
      n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, 
      n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, 
      n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, 
      n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, 
      n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, 
      n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, 
      n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, 
      n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, 
      n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, 
      n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, 
      n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, 
      n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, 
      n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, 
      n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, 
      n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, 
      n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, 
      n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, 
      n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, 
      n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, 
      n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, 
      n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, 
      n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, 
      n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, 
      n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, 
      n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, 
      n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, 
      n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, 
      n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, 
      n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, 
      n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, 
      n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, 
      n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, 
      n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, 
      n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, 
      n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, 
      n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, 
      n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, 
      n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, 
      n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, 
      n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, 
      n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, 
      n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, 
      n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, 
      n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, 
      n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, 
      n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, 
      n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, 
      n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, 
      n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, 
      n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, 
      n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, 
      n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, 
      n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, 
      n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, 
      n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, 
      n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, 
      n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, 
      n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, 
      n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, 
      n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, 
      n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, 
      n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, 
      n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, 
      n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, 
      n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, 
      n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, 
      n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, 
      n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, n_1792, 
      n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, 
      n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, 
      n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, 
      n_1820, n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828, 
      n_1829, n_1830, n_1831, n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, 
      n_1838, n_1839, n_1840, n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, 
      n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, 
      n_1856, n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, n_1863, n_1864, 
      n_1865, n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, 
      n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, 
      n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, 
      n_1892, n_1893, n_1894, n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, 
      n_1901, n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908, n_1909, 
      n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, 
      n_1919, n_1920, n_1921, n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, 
      n_1928, n_1929, n_1930, n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, 
      n_1937, n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, 
      n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, 
      n_1955, n_1956, n_1957, n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, 
      n_1964, n_1965, n_1966, n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, 
      n_1973, n_1974, n_1975, n_1976, n_1977, n_1978, n_1979, n_1980, n_1981, 
      n_1982, n_1983, n_1984, n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, 
      n_1991, n_1992, n_1993, n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, 
      n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, n_2007, n_2008, 
      n_2009, n_2010, n_2011, n_2012, n_2013, n_2014, n_2015, n_2016, n_2017, 
      n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, n_2024, n_2025, n_2026, 
      n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, 
      n_2036, n_2037, n_2038, n_2039, n_2040, n_2041, n_2042, n_2043, n_2044, 
      n_2045, n_2046, n_2047, n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, 
      n_2054, n_2055, n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, 
      n_2063, n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, 
      n_2072, n_2073, n_2074, n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, 
      n_2081, n_2082, n_2083, n_2084, n_2085, n_2086, n_2087, n_2088, n_2089, 
      n_2090, n_2091, n_2092, n_2093, n_2094, n_2095, n_2096, n_2097, n_2098, 
      n_2099, n_2100, n_2101, n_2102, n_2103, n_2104, n_2105, n_2106, n_2107, 
      n_2108, n_2109, n_2110, n_2111, n_2112, n_2113, n_2114, n_2115, n_2116, 
      n_2117, n_2118, n_2119, n_2120, n_2121, n_2122, n_2123, n_2124, n_2125, 
      n_2126, n_2127, n_2128, n_2129, n_2130, n_2131, n_2132, n_2133, n_2134, 
      n_2135, n_2136, n_2137, n_2138, n_2139, n_2140, n_2141, n_2142, n_2143, 
      n_2144, n_2145, n_2146, n_2147, n_2148, n_2149, n_2150, n_2151, n_2152, 
      n_2153, n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, n_2160, n_2161, 
      n_2162, n_2163, n_2164, n_2165, n_2166, n_2167, n_2168, n_2169, n_2170, 
      n_2171, n_2172, n_2173, n_2174, n_2175, n_2176, n_2177, n_2178, n_2179, 
      n_2180, n_2181, n_2182, n_2183, n_2184, n_2185, n_2186, n_2187, n_2188, 
      n_2189, n_2190, n_2191, n_2192, n_2193, n_2194, n_2195, n_2196, n_2197, 
      n_2198, n_2199, n_2200, n_2201, n_2202, n_2203, n_2204, n_2205, n_2206, 
      n_2207, n_2208, n_2209, n_2210, n_2211, n_2212, n_2213, n_2214, n_2215, 
      n_2216, n_2217, n_2218, n_2219, n_2220, n_2221, n_2222, n_2223, n_2224, 
      n_2225, n_2226, n_2227, n_2228, n_2229, n_2230, n_2231, n_2232, n_2233, 
      n_2234, n_2235, n_2236, n_2237, n_2238, n_2239, n_2240, n_2241, n_2242, 
      n_2243, n_2244, n_2245, n_2246, n_2247, n_2248, n_2249, n_2250, n_2251, 
      n_2252, n_2253, n_2254, n_2255, n_2256, n_2257, n_2258, n_2259, n_2260, 
      n_2261, n_2262, n_2263, n_2264, n_2265, n_2266, n_2267, n_2268, n_2269, 
      n_2270, n_2271, n_2272, n_2273, n_2274, n_2275, n_2276, n_2277, n_2278, 
      n_2279, n_2280, n_2281, n_2282, n_2283, n_2284, n_2285, n_2286, n_2287, 
      n_2288, n_2289, n_2290, n_2291, n_2292, n_2293, n_2294, n_2295, n_2296, 
      n_2297, n_2298, n_2299, n_2300, n_2301, n_2302, n_2303, n_2304, n_2305, 
      n_2306, n_2307, n_2308, n_2309, n_2310, n_2311, n_2312, n_2313, n_2314, 
      n_2315, n_2316, n_2317, n_2318, n_2319, n_2320, n_2321, n_2322, n_2323, 
      n_2324, n_2325, n_2326, n_2327, n_2328, n_2329, n_2330, n_2331, n_2332, 
      n_2333, n_2334, n_2335, n_2336, n_2337, n_2338, n_2339, n_2340, n_2341, 
      n_2342, n_2343, n_2344, n_2345, n_2346, n_2347, n_2348, n_2349, n_2350, 
      n_2351, n_2352, n_2353, n_2354, n_2355, n_2356, n_2357, n_2358, n_2359, 
      n_2360, n_2361, n_2362, n_2363, n_2364, n_2365, n_2366, n_2367, n_2368, 
      n_2369, n_2370, n_2371, n_2372, n_2373, n_2374, n_2375, n_2376, n_2377, 
      n_2378, n_2379, n_2380, n_2381, n_2382, n_2383, n_2384, n_2385, n_2386, 
      n_2387, n_2388, n_2389, n_2390, n_2391, n_2392, n_2393, n_2394, n_2395, 
      n_2396, n_2397, n_2398, n_2399, n_2400, n_2401, n_2402, n_2403, n_2404, 
      n_2405, n_2406, n_2407, n_2408, n_2409, n_2410, n_2411, n_2412, n_2413, 
      n_2414, n_2415, n_2416, n_2417, n_2418, n_2419, n_2420, n_2421, n_2422, 
      n_2423, n_2424, n_2425, n_2426, n_2427, n_2428, n_2429, n_2430, n_2431, 
      n_2432, n_2433, n_2434, n_2435, n_2436, n_2437, n_2438, n_2439, n_2440, 
      n_2441, n_2442, n_2443, n_2444, n_2445, n_2446, n_2447, n_2448, n_2449, 
      n_2450, n_2451, n_2452, n_2453, n_2454, n_2455, n_2456, n_2457, n_2458, 
      n_2459, n_2460, n_2461, n_2462, n_2463, n_2464, n_2465, n_2466, n_2467, 
      n_2468, n_2469, n_2470, n_2471, n_2472, n_2473, n_2474, n_2475, n_2476, 
      n_2477, n_2478, n_2479, n_2480, n_2481, n_2482, n_2483, n_2484, n_2485, 
      n_2486, n_2487, n_2488, n_2489, n_2490, n_2491, n_2492, n_2493, n_2494, 
      n_2495, n_2496, n_2497, n_2498, n_2499, n_2500, n_2501, n_2502, n_2503, 
      n_2504, n_2505, n_2506, n_2507, n_2508, n_2509, n_2510, n_2511, n_2512, 
      n_2513, n_2514, n_2515, n_2516, n_2517, n_2518, n_2519, n_2520, n_2521, 
      n_2522, n_2523, n_2524, n_2525, n_2526, n_2527, n_2528, n_2529, n_2530, 
      n_2531, n_2532, n_2533, n_2534, n_2535, n_2536, n_2537, n_2538, n_2539, 
      n_2540, n_2541, n_2542, n_2543, n_2544, n_2545, n_2546, n_2547, n_2548, 
      n_2549, n_2550, n_2551, n_2552, n_2553, n_2554, n_2555, n_2556, n_2557, 
      n_2558, n_2559, n_2560, n_2561, n_2562, n_2563, n_2564, n_2565, n_2566, 
      n_2567, n_2568, n_2569, n_2570, n_2571, n_2572, n_2573, n_2574, n_2575, 
      n_2576, n_2577, n_2578, n_2579, n_2580, n_2581, n_2582, n_2583, n_2584, 
      n_2585, n_2586, n_2587, n_2588, n_2589, n_2590, n_2591, n_2592, n_2593, 
      n_2594, n_2595, n_2596, n_2597, n_2598, n_2599, n_2600, n_2601, n_2602, 
      n_2603, n_2604, n_2605, n_2606, n_2607, n_2608, n_2609, n_2610, n_2611, 
      n_2612, n_2613, n_2614, n_2615, n_2616, n_2617, n_2618, n_2619, n_2620, 
      n_2621, n_2622, n_2623, n_2624, n_2625, n_2626, n_2627, n_2628, n_2629, 
      n_2630, n_2631, n_2632, n_2633, n_2634, n_2635, n_2636, n_2637, n_2638, 
      n_2639, n_2640, n_2641, n_2642, n_2643, n_2644, n_2645, n_2646, n_2647, 
      n_2648, n_2649, n_2650, n_2651, n_2652, n_2653, n_2654, n_2655, n_2656, 
      n_2657, n_2658, n_2659, n_2660, n_2661, n_2662, n_2663, n_2664, n_2665, 
      n_2666, n_2667, n_2668, n_2669, n_2670, n_2671, n_2672, n_2673, n_2674, 
      n_2675, n_2676, n_2677, n_2678, n_2679, n_2680, n_2681, n_2682, n_2683, 
      n_2684, n_2685, n_2686, n_2687, n_2688, n_2689, n_2690, n_2691, n_2692, 
      n_2693, n_2694, n_2695, n_2696, n_2697, n_2698, n_2699, n_2700, n_2701, 
      n_2702, n_2703, n_2704, n_2705, n_2706, n_2707, n_2708, n_2709, n_2710, 
      n_2711, n_2712, n_2713, n_2714, n_2715, n_2716, n_2717, n_2718, n_2719, 
      n_2720, n_2721, n_2722, n_2723, n_2724, n_2725, n_2726, n_2727, n_2728, 
      n_2729, n_2730, n_2731, n_2732, n_2733, n_2734, n_2735, n_2736, n_2737, 
      n_2738, n_2739, n_2740, n_2741, n_2742, n_2743, n_2744, n_2745, n_2746, 
      n_2747, n_2748, n_2749, n_2750, n_2751, n_2752, n_2753, n_2754, n_2755, 
      n_2756, n_2757, n_2758, n_2759, n_2760, n_2761, n_2762, n_2763, n_2764, 
      n_2765, n_2766, n_2767, n_2768, n_2769, n_2770, n_2771, n_2772, n_2773, 
      n_2774, n_2775, n_2776, n_2777, n_2778, n_2779, n_2780, n_2781, n_2782, 
      n_2783, n_2784, n_2785, n_2786, n_2787, n_2788, n_2789, n_2790, n_2791, 
      n_2792, n_2793, n_2794, n_2795, n_2796, n_2797, n_2798, n_2799, n_2800, 
      n_2801, n_2802, n_2803, n_2804, n_2805, n_2806, n_2807, n_2808, n_2809, 
      n_2810, n_2811, n_2812, n_2813, n_2814, n_2815, n_2816, n_2817, n_2818, 
      n_2819, n_2820, n_2821, n_2822, n_2823, n_2824, n_2825, n_2826, n_2827, 
      n_2828, n_2829, n_2830, n_2831, n_2832, n_2833, n_2834, n_2835, n_2836, 
      n_2837, n_2838, n_2839, n_2840, n_2841, n_2842, n_2843, n_2844, n_2845, 
      n_2846, n_2847, n_2848, n_2849, n_2850, n_2851, n_2852, n_2853, n_2854, 
      n_2855, n_2856, n_2857, n_2858, n_2859, n_2860, n_2861, n_2862, n_2863, 
      n_2864, n_2865, n_2866, n_2867, n_2868, n_2869, n_2870, n_2871, n_2872, 
      n_2873, n_2874, n_2875, n_2876, n_2877, n_2878, n_2879, n_2880, n_2881, 
      n_2882, n_2883, n_2884, n_2885, n_2886, n_2887, n_2888, n_2889, n_2890, 
      n_2891, n_2892, n_2893, n_2894, n_2895, n_2896, n_2897, n_2898, n_2899, 
      n_2900, n_2901, n_2902, n_2903, n_2904, n_2905, n_2906, n_2907, n_2908, 
      n_2909, n_2910, n_2911, n_2912, n_2913, n_2914, n_2915, n_2916, n_2917, 
      n_2918, n_2919, n_2920, n_2921, n_2922, n_2923, n_2924, n_2925, n_2926, 
      n_2927, n_2928, n_2929, n_2930, n_2931, n_2932, n_2933, n_2934, n_2935, 
      n_2936, n_2937, n_2938, n_2939, n_2940, n_2941, n_2942, n_2943, n_2944, 
      n_2945, n_2946, n_2947, n_2948, n_2949, n_2950, n_2951, n_2952, n_2953, 
      n_2954, n_2955, n_2956, n_2957, n_2958, n_2959, n_2960, n_2961, n_2962, 
      n_2963, n_2964, n_2965, n_2966, n_2967, n_2968, n_2969, n_2970, n_2971, 
      n_2972, n_2973, n_2974, n_2975, n_2976, n_2977, n_2978, n_2979, n_2980, 
      n_2981, n_2982, n_2983, n_2984, n_2985, n_2986, n_2987, n_2988, n_2989, 
      n_2990, n_2991, n_2992, n_2993, n_2994, n_2995, n_2996, n_2997, n_2998, 
      n_2999, n_3000, n_3001, n_3002, n_3003, n_3004, n_3005, n_3006, n_3007, 
      n_3008, n_3009, n_3010, n_3011, n_3012, n_3013, n_3014, n_3015, n_3016, 
      n_3017, n_3018, n_3019, n_3020, n_3021, n_3022, n_3023, n_3024, n_3025, 
      n_3026, n_3027, n_3028, n_3029, n_3030, n_3031, n_3032, n_3033, n_3034, 
      n_3035, n_3036, n_3037, n_3038, n_3039, n_3040, n_3041, n_3042, n_3043, 
      n_3044, n_3045, n_3046, n_3047, n_3048, n_3049, n_3050, n_3051, n_3052, 
      n_3053, n_3054, n_3055, n_3056, n_3057, n_3058, n_3059, n_3060, n_3061, 
      n_3062, n_3063, n_3064, n_3065, n_3066, n_3067, n_3068, n_3069, n_3070, 
      n_3071, n_3072, n_3073, n_3074, n_3075, n_3076, n_3077, n_3078, n_3079, 
      n_3080, n_3081, n_3082, n_3083, n_3084, n_3085, n_3086, n_3087, n_3088, 
      n_3089, n_3090, n_3091, n_3092, n_3093, n_3094, n_3095, n_3096, n_3097, 
      n_3098, n_3099, n_3100, n_3101, n_3102, n_3103, n_3104, n_3105, n_3106, 
      n_3107, n_3108, n_3109, n_3110, n_3111, n_3112, n_3113, n_3114, n_3115, 
      n_3116, n_3117, n_3118, n_3119, n_3120, n_3121, n_3122, n_3123, n_3124, 
      n_3125, n_3126, n_3127, n_3128, n_3129, n_3130, n_3131, n_3132, n_3133, 
      n_3134, n_3135, n_3136, n_3137, n_3138, n_3139, n_3140, n_3141, n_3142, 
      n_3143, n_3144, n_3145, n_3146, n_3147, n_3148, n_3149, n_3150, n_3151, 
      n_3152, n_3153, n_3154, n_3155 : std_logic;

begin
   
   i_BYTE_CNTR4_reg2 : FD1 port map( D => n6763, CP => CLK_I, Q => n1719, QN =>
                           n2505);
   i_BYTE_CNTR4_reg : FD1 port map( D => n6762, CP => CLK_I, Q => n1832, QN => 
                           n2506);
   FF_VALID_KEY_reg : FD1 port map( D => n4604, CP => CLK_I, Q => n_1000, QN =>
                           n4563);
   v_KEY32_IN_reg_31_inst : FD1 port map( D => n2421, CP => CLK_I, Q => 
                           v_KEY32_IN_31_port, QN => n_1001);
   v_KEY32_IN_reg_30_inst : FD1 port map( D => n2420, CP => CLK_I, Q => 
                           v_KEY32_IN_30_port, QN => n_1002);
   v_KEY32_IN_reg_29_inst : FD1 port map( D => n2419, CP => CLK_I, Q => 
                           v_KEY32_IN_29_port, QN => n_1003);
   v_KEY32_IN_reg_28_inst : FD1 port map( D => n2418, CP => CLK_I, Q => 
                           v_KEY32_IN_28_port, QN => n_1004);
   v_KEY32_IN_reg_27_inst : FD1 port map( D => n2417, CP => CLK_I, Q => 
                           v_KEY32_IN_27_port, QN => n_1005);
   v_KEY32_IN_reg_26_inst : FD1 port map( D => n2416, CP => CLK_I, Q => 
                           v_KEY32_IN_26_port, QN => n_1006);
   v_KEY32_IN_reg_25_inst : FD1 port map( D => n2415, CP => CLK_I, Q => 
                           v_KEY32_IN_25_port, QN => n_1007);
   v_KEY32_IN_reg_24_inst : FD1 port map( D => n2414, CP => CLK_I, Q => 
                           v_KEY32_IN_24_port, QN => n_1008);
   v_KEY32_IN_reg_23_inst : FD1 port map( D => n2429, CP => CLK_I, Q => 
                           v_KEY32_IN_23_port, QN => n_1009);
   v_KEY32_IN_reg_22_inst : FD1 port map( D => n2428, CP => CLK_I, Q => 
                           v_KEY32_IN_22_port, QN => n_1010);
   v_KEY32_IN_reg_21_inst : FD1 port map( D => n2427, CP => CLK_I, Q => 
                           v_KEY32_IN_21_port, QN => n_1011);
   v_KEY32_IN_reg_20_inst : FD1 port map( D => n2426, CP => CLK_I, Q => 
                           v_KEY32_IN_20_port, QN => n_1012);
   v_KEY32_IN_reg_19_inst : FD1 port map( D => n2425, CP => CLK_I, Q => 
                           v_KEY32_IN_19_port, QN => n_1013);
   v_KEY32_IN_reg_18_inst : FD1 port map( D => n2424, CP => CLK_I, Q => 
                           v_KEY32_IN_18_port, QN => n_1014);
   v_KEY32_IN_reg_17_inst : FD1 port map( D => n2423, CP => CLK_I, Q => 
                           v_KEY32_IN_17_port, QN => n_1015);
   v_KEY32_IN_reg_16_inst : FD1 port map( D => n2422, CP => CLK_I, Q => 
                           v_KEY32_IN_16_port, QN => n_1016);
   v_KEY32_IN_reg_15_inst : FD1 port map( D => n2438, CP => CLK_I, Q => 
                           v_KEY32_IN_15_port, QN => n_1017);
   v_KEY32_IN_reg_14_inst : FD1 port map( D => n2437, CP => CLK_I, Q => 
                           v_KEY32_IN_14_port, QN => n_1018);
   v_KEY32_IN_reg_13_inst : FD1 port map( D => n2436, CP => CLK_I, Q => 
                           v_KEY32_IN_13_port, QN => n_1019);
   v_KEY32_IN_reg_12_inst : FD1 port map( D => n2435, CP => CLK_I, Q => 
                           v_KEY32_IN_12_port, QN => n_1020);
   v_KEY32_IN_reg_11_inst : FD1 port map( D => n2434, CP => CLK_I, Q => 
                           v_KEY32_IN_11_port, QN => n_1021);
   v_KEY32_IN_reg_10_inst : FD1 port map( D => n2433, CP => CLK_I, Q => 
                           v_KEY32_IN_10_port, QN => n_1022);
   v_KEY32_IN_reg_9_inst : FD1 port map( D => n2432, CP => CLK_I, Q => 
                           v_KEY32_IN_9_port, QN => n_1023);
   v_KEY32_IN_reg_8_inst : FD1 port map( D => n2431, CP => CLK_I, Q => 
                           v_KEY32_IN_8_port, QN => n_1024);
   v_KEY32_IN_reg_7_inst : FD1 port map( D => n2413, CP => CLK_I, Q => 
                           v_KEY32_IN_7_port, QN => n_1025);
   v_KEY32_IN_reg_6_inst : FD1 port map( D => n2412, CP => CLK_I, Q => 
                           v_KEY32_IN_6_port, QN => n_1026);
   v_KEY32_IN_reg_5_inst : FD1 port map( D => n2411, CP => CLK_I, Q => 
                           v_KEY32_IN_5_port, QN => n_1027);
   v_KEY32_IN_reg_4_inst : FD1 port map( D => n2410, CP => CLK_I, Q => 
                           v_KEY32_IN_4_port, QN => n_1028);
   v_KEY32_IN_reg_3_inst : FD1 port map( D => n2409, CP => CLK_I, Q => 
                           v_KEY32_IN_3_port, QN => n_1029);
   v_KEY32_IN_reg_2_inst : FD1 port map( D => n2408, CP => CLK_I, Q => 
                           v_KEY32_IN_2_port, QN => n_1030);
   v_KEY32_IN_reg_1_inst : FD1 port map( D => n2407, CP => CLK_I, Q => 
                           v_KEY32_IN_1_port, QN => n_1031);
   v_KEY32_IN_reg_0_inst : FD1 port map( D => n2406, CP => CLK_I, Q => 
                           v_KEY32_IN_0_port, QN => n_1032);
   FF_GET_KEY_reg : FD1 port map( D => GET_KEY_I, CP => CLK_I, Q => n_1033, QN 
                           => n1793);
   v_SUB_WORD_reg_7_inst : FD1 port map( D => n4603, CP => CLK_I, Q => n_1034, 
                           QN => n2240);
   v_SUB_WORD_reg_6_inst : FD1 port map( D => n4602, CP => CLK_I, Q => n_1035, 
                           QN => n2183);
   v_SUB_WORD_reg_5_inst : FD1 port map( D => n4601, CP => CLK_I, Q => n_1036, 
                           QN => n2233);
   v_SUB_WORD_reg_4_inst : FD1 port map( D => n4600, CP => CLK_I, Q => n4561, 
                           QN => n2244);
   v_SUB_WORD_reg_3_inst : FD1 port map( D => n4599, CP => CLK_I, Q => n_1037, 
                           QN => n2220);
   v_SUB_WORD_reg_2_inst : FD1 port map( D => n4598, CP => CLK_I, Q => n_1038, 
                           QN => n2217);
   v_SUB_WORD_reg_1_inst : FD1 port map( D => n4597, CP => CLK_I, Q => n_1039, 
                           QN => n2205);
   v_SUB_WORD_reg_0_inst : FD1 port map( D => n4596, CP => CLK_I, Q => n_1040, 
                           QN => n2181);
   v_CALCULATION_CNTR_reg_0_inst : FD1 port map( D => n6665, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_0_port, QN => n2255);
   i_ROUND_reg : FD1 port map( D => n6729, CP => CLK_I, Q => n2091, QN => n6674
                           );
   START_CALCULATION_reg : FD1 port map( D => n6725, CP => CLK_I, Q => n_1041, 
                           QN => n6673);
   i_ROUND_reg4 : FD1 port map( D => n6728, CP => CLK_I, Q => n1833, QN => 
                           n6677);
   i_ROUND_reg3 : FD1 port map( D => n6727, CP => CLK_I, Q => n1875, QN => 
                           n6676);
   i_ROUND_reg2 : FD1 port map( D => n6726, CP => CLK_I, Q => n2050, QN => 
                           n6675);
   DONE_O_reg : FD1 port map( D => n6724, CP => CLK_I, Q => DONE_O, QN => n2507
                           );
   CALCULATION_reg : FD1 port map( D => n6723, CP => CLK_I, Q => n_1042, QN => 
                           n2031);
   v_CALCULATION_CNTR_reg_1_inst : FD1 port map( D => n6666, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_1_port, QN => n1882);
   v_CALCULATION_CNTR_reg_2_inst : FD1 port map( D => n6667, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_2_port, QN => n1877);
   v_CALCULATION_CNTR_reg_3_inst : FD1 port map( D => n6668, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_3_port, QN => n1883);
   v_CALCULATION_CNTR_reg_4_inst : FD1 port map( D => n6669, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_4_port, QN => n1844);
   v_CALCULATION_CNTR_reg_5_inst : FD1 port map( D => n2491, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_5_port, QN => n_1043);
   v_CALCULATION_CNTR_reg_6_inst : FD1 port map( D => n2492, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_6_port, QN => n2161);
   v_CALCULATION_CNTR_reg_7_inst : FD1 port map( D => n2494, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_7_port, QN => n_1044);
   i_INTERN_ADDR_RD0_reg6 : FD1 port map( D => n6722, CP => CLK_I, Q => 
                           i_INTERN_ADDR_RD05, QN => n6664);
   i_INTERN_ADDR_RD0_reg5 : FD1 port map( D => n6721, CP => CLK_I, Q => 
                           i_INTERN_ADDR_RD04, QN => n6663);
   i_INTERN_ADDR_RD0_reg4 : FD1 port map( D => n6720, CP => CLK_I, Q => 
                           i_INTERN_ADDR_RD03, QN => n6662);
   i_INTERN_ADDR_RD0_reg3 : FD1 port map( D => n6719, CP => CLK_I, Q => 
                           i_INTERN_ADDR_RD02, QN => n6661);
   i_INTERN_ADDR_RD0_reg2 : FD1 port map( D => n6718, CP => CLK_I, Q => 
                           i_INTERN_ADDR_RD01, QN => n6660);
   i_INTERN_ADDR_RD0_reg : FD1 port map( D => n6717, CP => CLK_I, Q => 
                           i_INTERN_ADDR_RD0, QN => n6659);
   SRAM_WREN0_reg : FD1 port map( D => n6716, CP => CLK_I, Q => n_1045, QN => 
                           n2509);
   i_SRAM_ADDR_WR0_reg : FD1 port map( D => n6715, CP => CLK_I, Q => 
                           i_SRAM_ADDR_WR0, QN => n6653);
   i_SRAM_ADDR_WR0_reg6 : FD1 port map( D => n6714, CP => CLK_I, Q => 
                           i_SRAM_ADDR_WR05, QN => n6658);
   i_SRAM_ADDR_WR0_reg5 : FD1 port map( D => n6713, CP => CLK_I, Q => 
                           i_SRAM_ADDR_WR04, QN => n6657);
   i_SRAM_ADDR_WR0_reg4 : FD1 port map( D => n6712, CP => CLK_I, Q => 
                           i_SRAM_ADDR_WR03, QN => n6656);
   i_SRAM_ADDR_WR0_reg3 : FD1 port map( D => n6711, CP => CLK_I, Q => 
                           i_SRAM_ADDR_WR02, QN => n6655);
   i_SRAM_ADDR_WR0_reg2 : FD1 port map( D => n6710, CP => CLK_I, Q => 
                           i_SRAM_ADDR_WR01, QN => n6654);
   v_TEMP_VECTOR_reg_7_inst : FD1 port map( D => n6702, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_7_port, QN => n_1046);
   KEY_EXPAN0_reg_63_7_inst : FD1 port map( D => n5116, CP => CLK_I, Q => 
                           n_1047, QN => n4519);
   KEY_EXPAN0_reg_62_7_inst : FD1 port map( D => n5115, CP => CLK_I, Q => 
                           n_1048, QN => n4518);
   KEY_EXPAN0_reg_61_7_inst : FD1 port map( D => n5114, CP => CLK_I, Q => 
                           n_1049, QN => n4521);
   KEY_EXPAN0_reg_60_7_inst : FD1 port map( D => n5113, CP => CLK_I, Q => 
                           n_1050, QN => n4520);
   KEY_EXPAN0_reg_59_7_inst : FD1 port map( D => n5112, CP => CLK_I, Q => 
                           n_1051, QN => n4523);
   KEY_EXPAN0_reg_58_7_inst : FD1 port map( D => n5111, CP => CLK_I, Q => 
                           n_1052, QN => n4522);
   KEY_EXPAN0_reg_57_7_inst : FD1 port map( D => n5110, CP => CLK_I, Q => 
                           n_1053, QN => n4525);
   KEY_EXPAN0_reg_56_7_inst : FD1 port map( D => n5109, CP => CLK_I, Q => 
                           n_1054, QN => n4524);
   KEY_EXPAN0_reg_55_7_inst : FD1 port map( D => n5108, CP => CLK_I, Q => 
                           n_1055, QN => n4511);
   KEY_EXPAN0_reg_54_7_inst : FD1 port map( D => n5107, CP => CLK_I, Q => 
                           n_1056, QN => n4510);
   KEY_EXPAN0_reg_53_7_inst : FD1 port map( D => n5106, CP => CLK_I, Q => 
                           n_1057, QN => n4513);
   KEY_EXPAN0_reg_52_7_inst : FD1 port map( D => n5105, CP => CLK_I, Q => 
                           n_1058, QN => n4512);
   KEY_EXPAN0_reg_51_7_inst : FD1 port map( D => n5104, CP => CLK_I, Q => 
                           n_1059, QN => n4515);
   KEY_EXPAN0_reg_50_7_inst : FD1 port map( D => n5103, CP => CLK_I, Q => 
                           n_1060, QN => n4514);
   KEY_EXPAN0_reg_49_7_inst : FD1 port map( D => n5102, CP => CLK_I, Q => 
                           n_1061, QN => n4517);
   KEY_EXPAN0_reg_48_7_inst : FD1 port map( D => n5101, CP => CLK_I, Q => 
                           n_1062, QN => n4516);
   KEY_EXPAN0_reg_47_7_inst : FD1 port map( D => n5100, CP => CLK_I, Q => 
                           n_1063, QN => n4503);
   KEY_EXPAN0_reg_46_7_inst : FD1 port map( D => n5099, CP => CLK_I, Q => 
                           n_1064, QN => n4502);
   KEY_EXPAN0_reg_45_7_inst : FD1 port map( D => n5098, CP => CLK_I, Q => 
                           n_1065, QN => n4505);
   KEY_EXPAN0_reg_44_7_inst : FD1 port map( D => n5097, CP => CLK_I, Q => 
                           n_1066, QN => n4504);
   KEY_EXPAN0_reg_43_7_inst : FD1 port map( D => n5096, CP => CLK_I, Q => 
                           n_1067, QN => n4507);
   KEY_EXPAN0_reg_42_7_inst : FD1 port map( D => n5095, CP => CLK_I, Q => 
                           n_1068, QN => n4506);
   KEY_EXPAN0_reg_41_7_inst : FD1 port map( D => n5094, CP => CLK_I, Q => 
                           n_1069, QN => n4509);
   KEY_EXPAN0_reg_40_7_inst : FD1 port map( D => n5093, CP => CLK_I, Q => 
                           n_1070, QN => n4508);
   KEY_EXPAN0_reg_39_7_inst : FD1 port map( D => n5092, CP => CLK_I, Q => 
                           n_1071, QN => n4495);
   KEY_EXPAN0_reg_38_7_inst : FD1 port map( D => n5091, CP => CLK_I, Q => 
                           n_1072, QN => n4494);
   KEY_EXPAN0_reg_37_7_inst : FD1 port map( D => n5090, CP => CLK_I, Q => 
                           n_1073, QN => n4497);
   KEY_EXPAN0_reg_36_7_inst : FD1 port map( D => n5089, CP => CLK_I, Q => 
                           n_1074, QN => n4496);
   KEY_EXPAN0_reg_35_7_inst : FD1 port map( D => n5088, CP => CLK_I, Q => 
                           n_1075, QN => n4499);
   KEY_EXPAN0_reg_34_7_inst : FD1 port map( D => n5087, CP => CLK_I, Q => 
                           n_1076, QN => n4498);
   KEY_EXPAN0_reg_33_7_inst : FD1 port map( D => n5086, CP => CLK_I, Q => 
                           n_1077, QN => n4501);
   KEY_EXPAN0_reg_32_7_inst : FD1 port map( D => n5085, CP => CLK_I, Q => 
                           n_1078, QN => n4500);
   KEY_EXPAN0_reg_31_7_inst : FD1 port map( D => n5084, CP => CLK_I, Q => 
                           n_1079, QN => n4551);
   KEY_EXPAN0_reg_30_7_inst : FD1 port map( D => n5083, CP => CLK_I, Q => 
                           n_1080, QN => n4550);
   KEY_EXPAN0_reg_29_7_inst : FD1 port map( D => n5082, CP => CLK_I, Q => 
                           n_1081, QN => n4553);
   KEY_EXPAN0_reg_28_7_inst : FD1 port map( D => n5081, CP => CLK_I, Q => 
                           n_1082, QN => n4552);
   KEY_EXPAN0_reg_27_7_inst : FD1 port map( D => n5080, CP => CLK_I, Q => 
                           n_1083, QN => n4555);
   KEY_EXPAN0_reg_26_7_inst : FD1 port map( D => n5079, CP => CLK_I, Q => 
                           n_1084, QN => n4554);
   KEY_EXPAN0_reg_25_7_inst : FD1 port map( D => n5078, CP => CLK_I, Q => 
                           n_1085, QN => n4557);
   KEY_EXPAN0_reg_24_7_inst : FD1 port map( D => n5077, CP => CLK_I, Q => 
                           n_1086, QN => n4556);
   KEY_EXPAN0_reg_23_7_inst : FD1 port map( D => n5076, CP => CLK_I, Q => 
                           n_1087, QN => n4543);
   KEY_EXPAN0_reg_22_7_inst : FD1 port map( D => n5075, CP => CLK_I, Q => 
                           n_1088, QN => n4542);
   KEY_EXPAN0_reg_21_7_inst : FD1 port map( D => n5074, CP => CLK_I, Q => 
                           n_1089, QN => n4545);
   KEY_EXPAN0_reg_20_7_inst : FD1 port map( D => n5073, CP => CLK_I, Q => 
                           n_1090, QN => n4544);
   KEY_EXPAN0_reg_19_7_inst : FD1 port map( D => n5072, CP => CLK_I, Q => 
                           n_1091, QN => n4547);
   KEY_EXPAN0_reg_18_7_inst : FD1 port map( D => n5071, CP => CLK_I, Q => 
                           n_1092, QN => n4546);
   KEY_EXPAN0_reg_17_7_inst : FD1 port map( D => n5070, CP => CLK_I, Q => 
                           n_1093, QN => n4549);
   KEY_EXPAN0_reg_16_7_inst : FD1 port map( D => n5069, CP => CLK_I, Q => 
                           n_1094, QN => n4548);
   KEY_EXPAN0_reg_15_7_inst : FD1 port map( D => n5068, CP => CLK_I, Q => 
                           n_1095, QN => n4535);
   KEY_EXPAN0_reg_14_7_inst : FD1 port map( D => n5067, CP => CLK_I, Q => 
                           n_1096, QN => n4534);
   KEY_EXPAN0_reg_13_7_inst : FD1 port map( D => n5066, CP => CLK_I, Q => 
                           n_1097, QN => n4537);
   KEY_EXPAN0_reg_12_7_inst : FD1 port map( D => n5065, CP => CLK_I, Q => 
                           n_1098, QN => n4536);
   KEY_EXPAN0_reg_11_7_inst : FD1 port map( D => n5064, CP => CLK_I, Q => 
                           n_1099, QN => n4539);
   KEY_EXPAN0_reg_10_7_inst : FD1 port map( D => n5063, CP => CLK_I, Q => 
                           n_1100, QN => n4538);
   KEY_EXPAN0_reg_9_7_inst : FD1 port map( D => n5062, CP => CLK_I, Q => n_1101
                           , QN => n4541);
   KEY_EXPAN0_reg_8_7_inst : FD1 port map( D => n5061, CP => CLK_I, Q => n_1102
                           , QN => n4540);
   KEY_EXPAN0_reg_7_7_inst : FD1 port map( D => n5060, CP => CLK_I, Q => n_1103
                           , QN => n4527);
   KEY_EXPAN0_reg_6_7_inst : FD1 port map( D => n5059, CP => CLK_I, Q => n_1104
                           , QN => n4526);
   KEY_EXPAN0_reg_5_7_inst : FD1 port map( D => n5058, CP => CLK_I, Q => n_1105
                           , QN => n4529);
   KEY_EXPAN0_reg_4_7_inst : FD1 port map( D => n5057, CP => CLK_I, Q => n_1106
                           , QN => n4528);
   KEY_EXPAN0_reg_3_7_inst : FD1 port map( D => n5056, CP => CLK_I, Q => n_1107
                           , QN => n4531);
   KEY_EXPAN0_reg_2_7_inst : FD1 port map( D => n5055, CP => CLK_I, Q => n_1108
                           , QN => n4530);
   KEY_EXPAN0_reg_1_7_inst : FD1 port map( D => n5054, CP => CLK_I, Q => n_1109
                           , QN => n4533);
   KEY_EXPAN0_reg_0_7_inst : FD1 port map( D => n5053, CP => CLK_I, Q => n_1110
                           , QN => n4532);
   v_KEY_COL_OUT0_reg_7_inst : FD1 port map( D => n4595, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_7_port, QN => n1866);
   v_TEMP_VECTOR_reg_31_inst : FD1 port map( D => n6678, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_31_port, QN => n_1111);
   KEY_EXPAN0_reg_63_31_inst : FD1 port map( D => n6652, CP => CLK_I, Q => 
                           n_1112, QN => n4455);
   KEY_EXPAN0_reg_62_31_inst : FD1 port map( D => n6651, CP => CLK_I, Q => 
                           n_1113, QN => n4454);
   KEY_EXPAN0_reg_61_31_inst : FD1 port map( D => n6650, CP => CLK_I, Q => 
                           n_1114, QN => n4457);
   KEY_EXPAN0_reg_60_31_inst : FD1 port map( D => n6649, CP => CLK_I, Q => 
                           n_1115, QN => n4456);
   KEY_EXPAN0_reg_59_31_inst : FD1 port map( D => n6648, CP => CLK_I, Q => 
                           n_1116, QN => n4459);
   KEY_EXPAN0_reg_58_31_inst : FD1 port map( D => n6647, CP => CLK_I, Q => 
                           n_1117, QN => n4458);
   KEY_EXPAN0_reg_57_31_inst : FD1 port map( D => n6646, CP => CLK_I, Q => 
                           n_1118, QN => n4461);
   KEY_EXPAN0_reg_56_31_inst : FD1 port map( D => n6645, CP => CLK_I, Q => 
                           n_1119, QN => n4460);
   KEY_EXPAN0_reg_55_31_inst : FD1 port map( D => n6644, CP => CLK_I, Q => 
                           n_1120, QN => n4447);
   KEY_EXPAN0_reg_54_31_inst : FD1 port map( D => n6643, CP => CLK_I, Q => 
                           n_1121, QN => n4446);
   KEY_EXPAN0_reg_53_31_inst : FD1 port map( D => n6642, CP => CLK_I, Q => 
                           n_1122, QN => n4449);
   KEY_EXPAN0_reg_52_31_inst : FD1 port map( D => n6641, CP => CLK_I, Q => 
                           n_1123, QN => n4448);
   KEY_EXPAN0_reg_51_31_inst : FD1 port map( D => n6640, CP => CLK_I, Q => 
                           n_1124, QN => n4451);
   KEY_EXPAN0_reg_50_31_inst : FD1 port map( D => n6639, CP => CLK_I, Q => 
                           n_1125, QN => n4450);
   KEY_EXPAN0_reg_49_31_inst : FD1 port map( D => n6638, CP => CLK_I, Q => 
                           n_1126, QN => n4453);
   KEY_EXPAN0_reg_48_31_inst : FD1 port map( D => n6637, CP => CLK_I, Q => 
                           n_1127, QN => n4452);
   KEY_EXPAN0_reg_47_31_inst : FD1 port map( D => n6636, CP => CLK_I, Q => 
                           n_1128, QN => n4439);
   KEY_EXPAN0_reg_46_31_inst : FD1 port map( D => n6635, CP => CLK_I, Q => 
                           n_1129, QN => n4438);
   KEY_EXPAN0_reg_45_31_inst : FD1 port map( D => n6634, CP => CLK_I, Q => 
                           n_1130, QN => n4441);
   KEY_EXPAN0_reg_44_31_inst : FD1 port map( D => n6633, CP => CLK_I, Q => 
                           n_1131, QN => n4440);
   KEY_EXPAN0_reg_43_31_inst : FD1 port map( D => n6632, CP => CLK_I, Q => 
                           n_1132, QN => n4443);
   KEY_EXPAN0_reg_42_31_inst : FD1 port map( D => n6631, CP => CLK_I, Q => 
                           n_1133, QN => n4442);
   KEY_EXPAN0_reg_41_31_inst : FD1 port map( D => n6630, CP => CLK_I, Q => 
                           n_1134, QN => n4445);
   KEY_EXPAN0_reg_40_31_inst : FD1 port map( D => n6629, CP => CLK_I, Q => 
                           n_1135, QN => n4444);
   KEY_EXPAN0_reg_39_31_inst : FD1 port map( D => n6628, CP => CLK_I, Q => 
                           n_1136, QN => n4431);
   KEY_EXPAN0_reg_38_31_inst : FD1 port map( D => n6627, CP => CLK_I, Q => 
                           n_1137, QN => n4430);
   KEY_EXPAN0_reg_37_31_inst : FD1 port map( D => n6626, CP => CLK_I, Q => 
                           n_1138, QN => n4433);
   KEY_EXPAN0_reg_36_31_inst : FD1 port map( D => n6625, CP => CLK_I, Q => 
                           n_1139, QN => n4432);
   KEY_EXPAN0_reg_35_31_inst : FD1 port map( D => n6624, CP => CLK_I, Q => 
                           n_1140, QN => n4435);
   KEY_EXPAN0_reg_34_31_inst : FD1 port map( D => n6623, CP => CLK_I, Q => 
                           n_1141, QN => n4434);
   KEY_EXPAN0_reg_33_31_inst : FD1 port map( D => n6622, CP => CLK_I, Q => 
                           n_1142, QN => n4437);
   KEY_EXPAN0_reg_32_31_inst : FD1 port map( D => n6621, CP => CLK_I, Q => 
                           n_1143, QN => n4436);
   KEY_EXPAN0_reg_31_31_inst : FD1 port map( D => n6620, CP => CLK_I, Q => 
                           n_1144, QN => n4487);
   KEY_EXPAN0_reg_30_31_inst : FD1 port map( D => n6619, CP => CLK_I, Q => 
                           n_1145, QN => n4486);
   KEY_EXPAN0_reg_29_31_inst : FD1 port map( D => n6618, CP => CLK_I, Q => 
                           n_1146, QN => n4489);
   KEY_EXPAN0_reg_28_31_inst : FD1 port map( D => n6617, CP => CLK_I, Q => 
                           n_1147, QN => n4488);
   KEY_EXPAN0_reg_27_31_inst : FD1 port map( D => n6616, CP => CLK_I, Q => 
                           n_1148, QN => n4491);
   KEY_EXPAN0_reg_26_31_inst : FD1 port map( D => n6615, CP => CLK_I, Q => 
                           n_1149, QN => n4490);
   KEY_EXPAN0_reg_25_31_inst : FD1 port map( D => n6614, CP => CLK_I, Q => 
                           n_1150, QN => n4493);
   KEY_EXPAN0_reg_24_31_inst : FD1 port map( D => n6613, CP => CLK_I, Q => 
                           n_1151, QN => n4492);
   KEY_EXPAN0_reg_23_31_inst : FD1 port map( D => n6612, CP => CLK_I, Q => 
                           n_1152, QN => n4479);
   KEY_EXPAN0_reg_22_31_inst : FD1 port map( D => n6611, CP => CLK_I, Q => 
                           n_1153, QN => n4478);
   KEY_EXPAN0_reg_21_31_inst : FD1 port map( D => n6610, CP => CLK_I, Q => 
                           n_1154, QN => n4481);
   KEY_EXPAN0_reg_20_31_inst : FD1 port map( D => n6609, CP => CLK_I, Q => 
                           n_1155, QN => n4480);
   KEY_EXPAN0_reg_19_31_inst : FD1 port map( D => n6608, CP => CLK_I, Q => 
                           n_1156, QN => n4483);
   KEY_EXPAN0_reg_18_31_inst : FD1 port map( D => n6607, CP => CLK_I, Q => 
                           n_1157, QN => n4482);
   KEY_EXPAN0_reg_17_31_inst : FD1 port map( D => n6606, CP => CLK_I, Q => 
                           n_1158, QN => n4485);
   KEY_EXPAN0_reg_16_31_inst : FD1 port map( D => n6605, CP => CLK_I, Q => 
                           n_1159, QN => n4484);
   KEY_EXPAN0_reg_15_31_inst : FD1 port map( D => n6604, CP => CLK_I, Q => 
                           n_1160, QN => n4471);
   KEY_EXPAN0_reg_14_31_inst : FD1 port map( D => n6603, CP => CLK_I, Q => 
                           n_1161, QN => n4470);
   KEY_EXPAN0_reg_13_31_inst : FD1 port map( D => n6602, CP => CLK_I, Q => 
                           n_1162, QN => n4473);
   KEY_EXPAN0_reg_12_31_inst : FD1 port map( D => n6601, CP => CLK_I, Q => 
                           n_1163, QN => n4472);
   KEY_EXPAN0_reg_11_31_inst : FD1 port map( D => n6600, CP => CLK_I, Q => 
                           n_1164, QN => n4475);
   KEY_EXPAN0_reg_10_31_inst : FD1 port map( D => n6599, CP => CLK_I, Q => 
                           n_1165, QN => n4474);
   KEY_EXPAN0_reg_9_31_inst : FD1 port map( D => n6598, CP => CLK_I, Q => 
                           n_1166, QN => n4477);
   KEY_EXPAN0_reg_8_31_inst : FD1 port map( D => n6597, CP => CLK_I, Q => 
                           n_1167, QN => n4476);
   KEY_EXPAN0_reg_7_31_inst : FD1 port map( D => n6596, CP => CLK_I, Q => 
                           n_1168, QN => n4463);
   KEY_EXPAN0_reg_6_31_inst : FD1 port map( D => n6595, CP => CLK_I, Q => 
                           n_1169, QN => n4462);
   KEY_EXPAN0_reg_5_31_inst : FD1 port map( D => n6594, CP => CLK_I, Q => 
                           n_1170, QN => n4465);
   KEY_EXPAN0_reg_4_31_inst : FD1 port map( D => n6593, CP => CLK_I, Q => 
                           n_1171, QN => n4464);
   KEY_EXPAN0_reg_3_31_inst : FD1 port map( D => n6592, CP => CLK_I, Q => 
                           n_1172, QN => n4467);
   KEY_EXPAN0_reg_2_31_inst : FD1 port map( D => n6591, CP => CLK_I, Q => 
                           n_1173, QN => n4466);
   KEY_EXPAN0_reg_1_31_inst : FD1 port map( D => n6590, CP => CLK_I, Q => 
                           n_1174, QN => n4469);
   KEY_EXPAN0_reg_0_31_inst : FD1 port map( D => n6589, CP => CLK_I, Q => 
                           n_1175, QN => n4468);
   v_KEY_COL_OUT0_reg_31_inst : FD1 port map( D => n4594, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_31_port, QN => n1941);
   v_TEMP_VECTOR_reg_23_inst : FD1 port map( D => n6686, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_23_port, QN => n_1176);
   KEY_EXPAN0_reg_63_23_inst : FD1 port map( D => n6140, CP => CLK_I, Q => 
                           n_1177, QN => n4391);
   KEY_EXPAN0_reg_62_23_inst : FD1 port map( D => n6139, CP => CLK_I, Q => 
                           n_1178, QN => n4390);
   KEY_EXPAN0_reg_61_23_inst : FD1 port map( D => n6138, CP => CLK_I, Q => 
                           n_1179, QN => n4393);
   KEY_EXPAN0_reg_60_23_inst : FD1 port map( D => n6137, CP => CLK_I, Q => 
                           n_1180, QN => n4392);
   KEY_EXPAN0_reg_59_23_inst : FD1 port map( D => n6136, CP => CLK_I, Q => 
                           n_1181, QN => n4395);
   KEY_EXPAN0_reg_58_23_inst : FD1 port map( D => n6135, CP => CLK_I, Q => 
                           n_1182, QN => n4394);
   KEY_EXPAN0_reg_57_23_inst : FD1 port map( D => n6134, CP => CLK_I, Q => 
                           n_1183, QN => n4397);
   KEY_EXPAN0_reg_56_23_inst : FD1 port map( D => n6133, CP => CLK_I, Q => 
                           n_1184, QN => n4396);
   KEY_EXPAN0_reg_55_23_inst : FD1 port map( D => n6132, CP => CLK_I, Q => 
                           n_1185, QN => n4383);
   KEY_EXPAN0_reg_54_23_inst : FD1 port map( D => n6131, CP => CLK_I, Q => 
                           n_1186, QN => n4382);
   KEY_EXPAN0_reg_53_23_inst : FD1 port map( D => n6130, CP => CLK_I, Q => 
                           n_1187, QN => n4385);
   KEY_EXPAN0_reg_52_23_inst : FD1 port map( D => n6129, CP => CLK_I, Q => 
                           n_1188, QN => n4384);
   KEY_EXPAN0_reg_51_23_inst : FD1 port map( D => n6128, CP => CLK_I, Q => 
                           n_1189, QN => n4387);
   KEY_EXPAN0_reg_50_23_inst : FD1 port map( D => n6127, CP => CLK_I, Q => 
                           n_1190, QN => n4386);
   KEY_EXPAN0_reg_49_23_inst : FD1 port map( D => n6126, CP => CLK_I, Q => 
                           n_1191, QN => n4389);
   KEY_EXPAN0_reg_48_23_inst : FD1 port map( D => n6125, CP => CLK_I, Q => 
                           n_1192, QN => n4388);
   KEY_EXPAN0_reg_47_23_inst : FD1 port map( D => n6124, CP => CLK_I, Q => 
                           n_1193, QN => n4375);
   KEY_EXPAN0_reg_46_23_inst : FD1 port map( D => n6123, CP => CLK_I, Q => 
                           n_1194, QN => n4374);
   KEY_EXPAN0_reg_45_23_inst : FD1 port map( D => n6122, CP => CLK_I, Q => 
                           n_1195, QN => n4377);
   KEY_EXPAN0_reg_44_23_inst : FD1 port map( D => n6121, CP => CLK_I, Q => 
                           n_1196, QN => n4376);
   KEY_EXPAN0_reg_43_23_inst : FD1 port map( D => n6120, CP => CLK_I, Q => 
                           n_1197, QN => n4379);
   KEY_EXPAN0_reg_42_23_inst : FD1 port map( D => n6119, CP => CLK_I, Q => 
                           n_1198, QN => n4378);
   KEY_EXPAN0_reg_41_23_inst : FD1 port map( D => n6118, CP => CLK_I, Q => 
                           n_1199, QN => n4381);
   KEY_EXPAN0_reg_40_23_inst : FD1 port map( D => n6117, CP => CLK_I, Q => 
                           n_1200, QN => n4380);
   KEY_EXPAN0_reg_39_23_inst : FD1 port map( D => n6116, CP => CLK_I, Q => 
                           n_1201, QN => n4367);
   KEY_EXPAN0_reg_38_23_inst : FD1 port map( D => n6115, CP => CLK_I, Q => 
                           n_1202, QN => n4366);
   KEY_EXPAN0_reg_37_23_inst : FD1 port map( D => n6114, CP => CLK_I, Q => 
                           n_1203, QN => n4369);
   KEY_EXPAN0_reg_36_23_inst : FD1 port map( D => n6113, CP => CLK_I, Q => 
                           n_1204, QN => n4368);
   KEY_EXPAN0_reg_35_23_inst : FD1 port map( D => n6112, CP => CLK_I, Q => 
                           n_1205, QN => n4371);
   KEY_EXPAN0_reg_34_23_inst : FD1 port map( D => n6111, CP => CLK_I, Q => 
                           n_1206, QN => n4370);
   KEY_EXPAN0_reg_33_23_inst : FD1 port map( D => n6110, CP => CLK_I, Q => 
                           n_1207, QN => n4373);
   KEY_EXPAN0_reg_32_23_inst : FD1 port map( D => n6109, CP => CLK_I, Q => 
                           n_1208, QN => n4372);
   KEY_EXPAN0_reg_31_23_inst : FD1 port map( D => n6108, CP => CLK_I, Q => 
                           n_1209, QN => n4423);
   KEY_EXPAN0_reg_30_23_inst : FD1 port map( D => n6107, CP => CLK_I, Q => 
                           n_1210, QN => n4422);
   KEY_EXPAN0_reg_29_23_inst : FD1 port map( D => n6106, CP => CLK_I, Q => 
                           n_1211, QN => n4425);
   KEY_EXPAN0_reg_28_23_inst : FD1 port map( D => n6105, CP => CLK_I, Q => 
                           n_1212, QN => n4424);
   KEY_EXPAN0_reg_27_23_inst : FD1 port map( D => n6104, CP => CLK_I, Q => 
                           n_1213, QN => n4427);
   KEY_EXPAN0_reg_26_23_inst : FD1 port map( D => n6103, CP => CLK_I, Q => 
                           n_1214, QN => n4426);
   KEY_EXPAN0_reg_25_23_inst : FD1 port map( D => n6102, CP => CLK_I, Q => 
                           n_1215, QN => n4429);
   KEY_EXPAN0_reg_24_23_inst : FD1 port map( D => n6101, CP => CLK_I, Q => 
                           n_1216, QN => n4428);
   KEY_EXPAN0_reg_23_23_inst : FD1 port map( D => n6100, CP => CLK_I, Q => 
                           n_1217, QN => n4415);
   KEY_EXPAN0_reg_22_23_inst : FD1 port map( D => n6099, CP => CLK_I, Q => 
                           n_1218, QN => n4414);
   KEY_EXPAN0_reg_21_23_inst : FD1 port map( D => n6098, CP => CLK_I, Q => 
                           n_1219, QN => n4417);
   KEY_EXPAN0_reg_20_23_inst : FD1 port map( D => n6097, CP => CLK_I, Q => 
                           n_1220, QN => n4416);
   KEY_EXPAN0_reg_19_23_inst : FD1 port map( D => n6096, CP => CLK_I, Q => 
                           n_1221, QN => n4419);
   KEY_EXPAN0_reg_18_23_inst : FD1 port map( D => n6095, CP => CLK_I, Q => 
                           n_1222, QN => n4418);
   KEY_EXPAN0_reg_17_23_inst : FD1 port map( D => n6094, CP => CLK_I, Q => 
                           n_1223, QN => n4421);
   KEY_EXPAN0_reg_16_23_inst : FD1 port map( D => n6093, CP => CLK_I, Q => 
                           n_1224, QN => n4420);
   KEY_EXPAN0_reg_15_23_inst : FD1 port map( D => n6092, CP => CLK_I, Q => 
                           n_1225, QN => n4407);
   KEY_EXPAN0_reg_14_23_inst : FD1 port map( D => n6091, CP => CLK_I, Q => 
                           n_1226, QN => n4406);
   KEY_EXPAN0_reg_13_23_inst : FD1 port map( D => n6090, CP => CLK_I, Q => 
                           n_1227, QN => n4409);
   KEY_EXPAN0_reg_12_23_inst : FD1 port map( D => n6089, CP => CLK_I, Q => 
                           n_1228, QN => n4408);
   KEY_EXPAN0_reg_11_23_inst : FD1 port map( D => n6088, CP => CLK_I, Q => 
                           n_1229, QN => n4411);
   KEY_EXPAN0_reg_10_23_inst : FD1 port map( D => n6087, CP => CLK_I, Q => 
                           n_1230, QN => n4410);
   KEY_EXPAN0_reg_9_23_inst : FD1 port map( D => n6086, CP => CLK_I, Q => 
                           n_1231, QN => n4413);
   KEY_EXPAN0_reg_8_23_inst : FD1 port map( D => n6085, CP => CLK_I, Q => 
                           n_1232, QN => n4412);
   KEY_EXPAN0_reg_7_23_inst : FD1 port map( D => n6084, CP => CLK_I, Q => 
                           n_1233, QN => n4399);
   KEY_EXPAN0_reg_6_23_inst : FD1 port map( D => n6083, CP => CLK_I, Q => 
                           n_1234, QN => n4398);
   KEY_EXPAN0_reg_5_23_inst : FD1 port map( D => n6082, CP => CLK_I, Q => 
                           n_1235, QN => n4401);
   KEY_EXPAN0_reg_4_23_inst : FD1 port map( D => n6081, CP => CLK_I, Q => 
                           n_1236, QN => n4400);
   KEY_EXPAN0_reg_3_23_inst : FD1 port map( D => n6080, CP => CLK_I, Q => 
                           n_1237, QN => n4403);
   KEY_EXPAN0_reg_2_23_inst : FD1 port map( D => n6079, CP => CLK_I, Q => 
                           n_1238, QN => n4402);
   KEY_EXPAN0_reg_1_23_inst : FD1 port map( D => n6078, CP => CLK_I, Q => 
                           n_1239, QN => n4405);
   KEY_EXPAN0_reg_0_23_inst : FD1 port map( D => n6077, CP => CLK_I, Q => 
                           n_1240, QN => n4404);
   v_KEY_COL_OUT0_reg_23_inst : FD1 port map( D => n4593, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_23_port, QN => n1917);
   v_TEMP_VECTOR_reg_15_inst : FD1 port map( D => n6694, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_15_port, QN => n_1241);
   KEY_EXPAN0_reg_63_15_inst : FD1 port map( D => n5628, CP => CLK_I, Q => 
                           n_1242, QN => n4327);
   KEY_EXPAN0_reg_62_15_inst : FD1 port map( D => n5627, CP => CLK_I, Q => 
                           n_1243, QN => n4326);
   KEY_EXPAN0_reg_61_15_inst : FD1 port map( D => n5626, CP => CLK_I, Q => 
                           n_1244, QN => n4329);
   KEY_EXPAN0_reg_60_15_inst : FD1 port map( D => n5625, CP => CLK_I, Q => 
                           n_1245, QN => n4328);
   KEY_EXPAN0_reg_59_15_inst : FD1 port map( D => n5624, CP => CLK_I, Q => 
                           n_1246, QN => n4331);
   KEY_EXPAN0_reg_58_15_inst : FD1 port map( D => n5623, CP => CLK_I, Q => 
                           n_1247, QN => n4330);
   KEY_EXPAN0_reg_57_15_inst : FD1 port map( D => n5622, CP => CLK_I, Q => 
                           n_1248, QN => n4333);
   KEY_EXPAN0_reg_56_15_inst : FD1 port map( D => n5621, CP => CLK_I, Q => 
                           n_1249, QN => n4332);
   KEY_EXPAN0_reg_55_15_inst : FD1 port map( D => n5620, CP => CLK_I, Q => 
                           n_1250, QN => n4319);
   KEY_EXPAN0_reg_54_15_inst : FD1 port map( D => n5619, CP => CLK_I, Q => 
                           n_1251, QN => n4318);
   KEY_EXPAN0_reg_53_15_inst : FD1 port map( D => n5618, CP => CLK_I, Q => 
                           n_1252, QN => n4321);
   KEY_EXPAN0_reg_52_15_inst : FD1 port map( D => n5617, CP => CLK_I, Q => 
                           n_1253, QN => n4320);
   KEY_EXPAN0_reg_51_15_inst : FD1 port map( D => n5616, CP => CLK_I, Q => 
                           n_1254, QN => n4323);
   KEY_EXPAN0_reg_50_15_inst : FD1 port map( D => n5615, CP => CLK_I, Q => 
                           n_1255, QN => n4322);
   KEY_EXPAN0_reg_49_15_inst : FD1 port map( D => n5614, CP => CLK_I, Q => 
                           n_1256, QN => n4325);
   KEY_EXPAN0_reg_48_15_inst : FD1 port map( D => n5613, CP => CLK_I, Q => 
                           n_1257, QN => n4324);
   KEY_EXPAN0_reg_47_15_inst : FD1 port map( D => n5612, CP => CLK_I, Q => 
                           n_1258, QN => n4311);
   KEY_EXPAN0_reg_46_15_inst : FD1 port map( D => n5611, CP => CLK_I, Q => 
                           n_1259, QN => n4310);
   KEY_EXPAN0_reg_45_15_inst : FD1 port map( D => n5610, CP => CLK_I, Q => 
                           n_1260, QN => n4313);
   KEY_EXPAN0_reg_44_15_inst : FD1 port map( D => n5609, CP => CLK_I, Q => 
                           n_1261, QN => n4312);
   KEY_EXPAN0_reg_43_15_inst : FD1 port map( D => n5608, CP => CLK_I, Q => 
                           n_1262, QN => n4315);
   KEY_EXPAN0_reg_42_15_inst : FD1 port map( D => n5607, CP => CLK_I, Q => 
                           n_1263, QN => n4314);
   KEY_EXPAN0_reg_41_15_inst : FD1 port map( D => n5606, CP => CLK_I, Q => 
                           n_1264, QN => n4317);
   KEY_EXPAN0_reg_40_15_inst : FD1 port map( D => n5605, CP => CLK_I, Q => 
                           n_1265, QN => n4316);
   KEY_EXPAN0_reg_39_15_inst : FD1 port map( D => n5604, CP => CLK_I, Q => 
                           n_1266, QN => n4303);
   KEY_EXPAN0_reg_38_15_inst : FD1 port map( D => n5603, CP => CLK_I, Q => 
                           n_1267, QN => n4302);
   KEY_EXPAN0_reg_37_15_inst : FD1 port map( D => n5602, CP => CLK_I, Q => 
                           n_1268, QN => n4305);
   KEY_EXPAN0_reg_36_15_inst : FD1 port map( D => n5601, CP => CLK_I, Q => 
                           n_1269, QN => n4304);
   KEY_EXPAN0_reg_35_15_inst : FD1 port map( D => n5600, CP => CLK_I, Q => 
                           n_1270, QN => n4307);
   KEY_EXPAN0_reg_34_15_inst : FD1 port map( D => n5599, CP => CLK_I, Q => 
                           n_1271, QN => n4306);
   KEY_EXPAN0_reg_33_15_inst : FD1 port map( D => n5598, CP => CLK_I, Q => 
                           n_1272, QN => n4309);
   KEY_EXPAN0_reg_32_15_inst : FD1 port map( D => n5597, CP => CLK_I, Q => 
                           n_1273, QN => n4308);
   KEY_EXPAN0_reg_31_15_inst : FD1 port map( D => n5596, CP => CLK_I, Q => 
                           n_1274, QN => n4359);
   KEY_EXPAN0_reg_30_15_inst : FD1 port map( D => n5595, CP => CLK_I, Q => 
                           n_1275, QN => n4358);
   KEY_EXPAN0_reg_29_15_inst : FD1 port map( D => n5594, CP => CLK_I, Q => 
                           n_1276, QN => n4361);
   KEY_EXPAN0_reg_28_15_inst : FD1 port map( D => n5593, CP => CLK_I, Q => 
                           n_1277, QN => n4360);
   KEY_EXPAN0_reg_27_15_inst : FD1 port map( D => n5592, CP => CLK_I, Q => 
                           n_1278, QN => n4363);
   KEY_EXPAN0_reg_26_15_inst : FD1 port map( D => n5591, CP => CLK_I, Q => 
                           n_1279, QN => n4362);
   KEY_EXPAN0_reg_25_15_inst : FD1 port map( D => n5590, CP => CLK_I, Q => 
                           n_1280, QN => n4365);
   KEY_EXPAN0_reg_24_15_inst : FD1 port map( D => n5589, CP => CLK_I, Q => 
                           n_1281, QN => n4364);
   KEY_EXPAN0_reg_23_15_inst : FD1 port map( D => n5588, CP => CLK_I, Q => 
                           n_1282, QN => n4351);
   KEY_EXPAN0_reg_22_15_inst : FD1 port map( D => n5587, CP => CLK_I, Q => 
                           n_1283, QN => n4350);
   KEY_EXPAN0_reg_21_15_inst : FD1 port map( D => n5586, CP => CLK_I, Q => 
                           n_1284, QN => n4353);
   KEY_EXPAN0_reg_20_15_inst : FD1 port map( D => n5585, CP => CLK_I, Q => 
                           n_1285, QN => n4352);
   KEY_EXPAN0_reg_19_15_inst : FD1 port map( D => n5584, CP => CLK_I, Q => 
                           n_1286, QN => n4355);
   KEY_EXPAN0_reg_18_15_inst : FD1 port map( D => n5583, CP => CLK_I, Q => 
                           n_1287, QN => n4354);
   KEY_EXPAN0_reg_17_15_inst : FD1 port map( D => n5582, CP => CLK_I, Q => 
                           n_1288, QN => n4357);
   KEY_EXPAN0_reg_16_15_inst : FD1 port map( D => n5581, CP => CLK_I, Q => 
                           n_1289, QN => n4356);
   KEY_EXPAN0_reg_15_15_inst : FD1 port map( D => n5580, CP => CLK_I, Q => 
                           n_1290, QN => n4343);
   KEY_EXPAN0_reg_14_15_inst : FD1 port map( D => n5579, CP => CLK_I, Q => 
                           n_1291, QN => n4342);
   KEY_EXPAN0_reg_13_15_inst : FD1 port map( D => n5578, CP => CLK_I, Q => 
                           n_1292, QN => n4345);
   KEY_EXPAN0_reg_12_15_inst : FD1 port map( D => n5577, CP => CLK_I, Q => 
                           n_1293, QN => n4344);
   KEY_EXPAN0_reg_11_15_inst : FD1 port map( D => n5576, CP => CLK_I, Q => 
                           n_1294, QN => n4347);
   KEY_EXPAN0_reg_10_15_inst : FD1 port map( D => n5575, CP => CLK_I, Q => 
                           n_1295, QN => n4346);
   KEY_EXPAN0_reg_9_15_inst : FD1 port map( D => n5574, CP => CLK_I, Q => 
                           n_1296, QN => n4349);
   KEY_EXPAN0_reg_8_15_inst : FD1 port map( D => n5573, CP => CLK_I, Q => 
                           n_1297, QN => n4348);
   KEY_EXPAN0_reg_7_15_inst : FD1 port map( D => n5572, CP => CLK_I, Q => 
                           n_1298, QN => n4335);
   KEY_EXPAN0_reg_6_15_inst : FD1 port map( D => n5571, CP => CLK_I, Q => 
                           n_1299, QN => n4334);
   KEY_EXPAN0_reg_5_15_inst : FD1 port map( D => n5570, CP => CLK_I, Q => 
                           n_1300, QN => n4337);
   KEY_EXPAN0_reg_4_15_inst : FD1 port map( D => n5569, CP => CLK_I, Q => 
                           n_1301, QN => n4336);
   KEY_EXPAN0_reg_3_15_inst : FD1 port map( D => n5568, CP => CLK_I, Q => 
                           n_1302, QN => n4339);
   KEY_EXPAN0_reg_2_15_inst : FD1 port map( D => n5567, CP => CLK_I, Q => 
                           n_1303, QN => n4338);
   KEY_EXPAN0_reg_1_15_inst : FD1 port map( D => n5566, CP => CLK_I, Q => 
                           n_1304, QN => n4341);
   KEY_EXPAN0_reg_0_15_inst : FD1 port map( D => n5565, CP => CLK_I, Q => 
                           n_1305, QN => n4340);
   v_KEY_COL_OUT0_reg_15_inst : FD1 port map( D => n4592, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_15_port, QN => n1908);
   v_TEMP_VECTOR_reg_6_inst : FD1 port map( D => n6703, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_6_port, QN => n2121);
   KEY_EXPAN0_reg_63_6_inst : FD1 port map( D => n5052, CP => CLK_I, Q => 
                           n_1306, QN => n4263);
   KEY_EXPAN0_reg_62_6_inst : FD1 port map( D => n5051, CP => CLK_I, Q => 
                           n_1307, QN => n4262);
   KEY_EXPAN0_reg_61_6_inst : FD1 port map( D => n5050, CP => CLK_I, Q => 
                           n_1308, QN => n4265);
   KEY_EXPAN0_reg_60_6_inst : FD1 port map( D => n5049, CP => CLK_I, Q => 
                           n_1309, QN => n4264);
   KEY_EXPAN0_reg_59_6_inst : FD1 port map( D => n5048, CP => CLK_I, Q => 
                           n_1310, QN => n4267);
   KEY_EXPAN0_reg_58_6_inst : FD1 port map( D => n5047, CP => CLK_I, Q => 
                           n_1311, QN => n4266);
   KEY_EXPAN0_reg_57_6_inst : FD1 port map( D => n5046, CP => CLK_I, Q => 
                           n_1312, QN => n4269);
   KEY_EXPAN0_reg_56_6_inst : FD1 port map( D => n5045, CP => CLK_I, Q => 
                           n_1313, QN => n4268);
   KEY_EXPAN0_reg_55_6_inst : FD1 port map( D => n5044, CP => CLK_I, Q => 
                           n_1314, QN => n4255);
   KEY_EXPAN0_reg_54_6_inst : FD1 port map( D => n5043, CP => CLK_I, Q => 
                           n_1315, QN => n4254);
   KEY_EXPAN0_reg_53_6_inst : FD1 port map( D => n5042, CP => CLK_I, Q => 
                           n_1316, QN => n4257);
   KEY_EXPAN0_reg_52_6_inst : FD1 port map( D => n5041, CP => CLK_I, Q => 
                           n_1317, QN => n4256);
   KEY_EXPAN0_reg_51_6_inst : FD1 port map( D => n5040, CP => CLK_I, Q => 
                           n_1318, QN => n4259);
   KEY_EXPAN0_reg_50_6_inst : FD1 port map( D => n5039, CP => CLK_I, Q => 
                           n_1319, QN => n4258);
   KEY_EXPAN0_reg_49_6_inst : FD1 port map( D => n5038, CP => CLK_I, Q => 
                           n_1320, QN => n4261);
   KEY_EXPAN0_reg_48_6_inst : FD1 port map( D => n5037, CP => CLK_I, Q => 
                           n_1321, QN => n4260);
   KEY_EXPAN0_reg_47_6_inst : FD1 port map( D => n5036, CP => CLK_I, Q => 
                           n_1322, QN => n4247);
   KEY_EXPAN0_reg_46_6_inst : FD1 port map( D => n5035, CP => CLK_I, Q => 
                           n_1323, QN => n4246);
   KEY_EXPAN0_reg_45_6_inst : FD1 port map( D => n5034, CP => CLK_I, Q => 
                           n_1324, QN => n4249);
   KEY_EXPAN0_reg_44_6_inst : FD1 port map( D => n5033, CP => CLK_I, Q => 
                           n_1325, QN => n4248);
   KEY_EXPAN0_reg_43_6_inst : FD1 port map( D => n5032, CP => CLK_I, Q => 
                           n_1326, QN => n4251);
   KEY_EXPAN0_reg_42_6_inst : FD1 port map( D => n5031, CP => CLK_I, Q => 
                           n_1327, QN => n4250);
   KEY_EXPAN0_reg_41_6_inst : FD1 port map( D => n5030, CP => CLK_I, Q => 
                           n_1328, QN => n4253);
   KEY_EXPAN0_reg_40_6_inst : FD1 port map( D => n5029, CP => CLK_I, Q => 
                           n_1329, QN => n4252);
   KEY_EXPAN0_reg_39_6_inst : FD1 port map( D => n5028, CP => CLK_I, Q => 
                           n_1330, QN => n4239);
   KEY_EXPAN0_reg_38_6_inst : FD1 port map( D => n5027, CP => CLK_I, Q => 
                           n_1331, QN => n4238);
   KEY_EXPAN0_reg_37_6_inst : FD1 port map( D => n5026, CP => CLK_I, Q => 
                           n_1332, QN => n4241);
   KEY_EXPAN0_reg_36_6_inst : FD1 port map( D => n5025, CP => CLK_I, Q => 
                           n_1333, QN => n4240);
   KEY_EXPAN0_reg_35_6_inst : FD1 port map( D => n5024, CP => CLK_I, Q => 
                           n_1334, QN => n4243);
   KEY_EXPAN0_reg_34_6_inst : FD1 port map( D => n5023, CP => CLK_I, Q => 
                           n_1335, QN => n4242);
   KEY_EXPAN0_reg_33_6_inst : FD1 port map( D => n5022, CP => CLK_I, Q => 
                           n_1336, QN => n4245);
   KEY_EXPAN0_reg_32_6_inst : FD1 port map( D => n5021, CP => CLK_I, Q => 
                           n_1337, QN => n4244);
   KEY_EXPAN0_reg_31_6_inst : FD1 port map( D => n5020, CP => CLK_I, Q => 
                           n_1338, QN => n4295);
   KEY_EXPAN0_reg_30_6_inst : FD1 port map( D => n5019, CP => CLK_I, Q => 
                           n_1339, QN => n4294);
   KEY_EXPAN0_reg_29_6_inst : FD1 port map( D => n5018, CP => CLK_I, Q => 
                           n_1340, QN => n4297);
   KEY_EXPAN0_reg_28_6_inst : FD1 port map( D => n5017, CP => CLK_I, Q => 
                           n_1341, QN => n4296);
   KEY_EXPAN0_reg_27_6_inst : FD1 port map( D => n5016, CP => CLK_I, Q => 
                           n_1342, QN => n4299);
   KEY_EXPAN0_reg_26_6_inst : FD1 port map( D => n5015, CP => CLK_I, Q => 
                           n_1343, QN => n4298);
   KEY_EXPAN0_reg_25_6_inst : FD1 port map( D => n5014, CP => CLK_I, Q => 
                           n_1344, QN => n4301);
   KEY_EXPAN0_reg_24_6_inst : FD1 port map( D => n5013, CP => CLK_I, Q => 
                           n_1345, QN => n4300);
   KEY_EXPAN0_reg_23_6_inst : FD1 port map( D => n5012, CP => CLK_I, Q => 
                           n_1346, QN => n4287);
   KEY_EXPAN0_reg_22_6_inst : FD1 port map( D => n5011, CP => CLK_I, Q => 
                           n_1347, QN => n4286);
   KEY_EXPAN0_reg_21_6_inst : FD1 port map( D => n5010, CP => CLK_I, Q => 
                           n_1348, QN => n4289);
   KEY_EXPAN0_reg_20_6_inst : FD1 port map( D => n5009, CP => CLK_I, Q => 
                           n_1349, QN => n4288);
   KEY_EXPAN0_reg_19_6_inst : FD1 port map( D => n5008, CP => CLK_I, Q => 
                           n_1350, QN => n4291);
   KEY_EXPAN0_reg_18_6_inst : FD1 port map( D => n5007, CP => CLK_I, Q => 
                           n_1351, QN => n4290);
   KEY_EXPAN0_reg_17_6_inst : FD1 port map( D => n5006, CP => CLK_I, Q => 
                           n_1352, QN => n4293);
   KEY_EXPAN0_reg_16_6_inst : FD1 port map( D => n5005, CP => CLK_I, Q => 
                           n_1353, QN => n4292);
   KEY_EXPAN0_reg_15_6_inst : FD1 port map( D => n5004, CP => CLK_I, Q => 
                           n_1354, QN => n4279);
   KEY_EXPAN0_reg_14_6_inst : FD1 port map( D => n5003, CP => CLK_I, Q => 
                           n_1355, QN => n4278);
   KEY_EXPAN0_reg_13_6_inst : FD1 port map( D => n5002, CP => CLK_I, Q => 
                           n_1356, QN => n4281);
   KEY_EXPAN0_reg_12_6_inst : FD1 port map( D => n5001, CP => CLK_I, Q => 
                           n_1357, QN => n4280);
   KEY_EXPAN0_reg_11_6_inst : FD1 port map( D => n5000, CP => CLK_I, Q => 
                           n_1358, QN => n4283);
   KEY_EXPAN0_reg_10_6_inst : FD1 port map( D => n4999, CP => CLK_I, Q => 
                           n_1359, QN => n4282);
   KEY_EXPAN0_reg_9_6_inst : FD1 port map( D => n4998, CP => CLK_I, Q => n_1360
                           , QN => n4285);
   KEY_EXPAN0_reg_8_6_inst : FD1 port map( D => n4997, CP => CLK_I, Q => n_1361
                           , QN => n4284);
   KEY_EXPAN0_reg_7_6_inst : FD1 port map( D => n4996, CP => CLK_I, Q => n_1362
                           , QN => n4271);
   KEY_EXPAN0_reg_6_6_inst : FD1 port map( D => n4995, CP => CLK_I, Q => n_1363
                           , QN => n4270);
   KEY_EXPAN0_reg_5_6_inst : FD1 port map( D => n4994, CP => CLK_I, Q => n_1364
                           , QN => n4273);
   KEY_EXPAN0_reg_4_6_inst : FD1 port map( D => n4993, CP => CLK_I, Q => n_1365
                           , QN => n4272);
   KEY_EXPAN0_reg_3_6_inst : FD1 port map( D => n4992, CP => CLK_I, Q => n_1366
                           , QN => n4275);
   KEY_EXPAN0_reg_2_6_inst : FD1 port map( D => n4991, CP => CLK_I, Q => n_1367
                           , QN => n4274);
   KEY_EXPAN0_reg_1_6_inst : FD1 port map( D => n4990, CP => CLK_I, Q => n_1368
                           , QN => n4277);
   KEY_EXPAN0_reg_0_6_inst : FD1 port map( D => n4989, CP => CLK_I, Q => n_1369
                           , QN => n4276);
   v_KEY_COL_OUT0_reg_6_inst : FD1 port map( D => n4591, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_6_port, QN => n1861);
   v_TEMP_VECTOR_reg_30_inst : FD1 port map( D => n6679, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_30_port, QN => n_1370);
   KEY_EXPAN0_reg_63_30_inst : FD1 port map( D => n6588, CP => CLK_I, Q => 
                           n_1371, QN => n4199);
   KEY_EXPAN0_reg_62_30_inst : FD1 port map( D => n6587, CP => CLK_I, Q => 
                           n_1372, QN => n4198);
   KEY_EXPAN0_reg_61_30_inst : FD1 port map( D => n6586, CP => CLK_I, Q => 
                           n_1373, QN => n4201);
   KEY_EXPAN0_reg_60_30_inst : FD1 port map( D => n6585, CP => CLK_I, Q => 
                           n_1374, QN => n4200);
   KEY_EXPAN0_reg_59_30_inst : FD1 port map( D => n6584, CP => CLK_I, Q => 
                           n_1375, QN => n4203);
   KEY_EXPAN0_reg_58_30_inst : FD1 port map( D => n6583, CP => CLK_I, Q => 
                           n_1376, QN => n4202);
   KEY_EXPAN0_reg_57_30_inst : FD1 port map( D => n6582, CP => CLK_I, Q => 
                           n_1377, QN => n4205);
   KEY_EXPAN0_reg_56_30_inst : FD1 port map( D => n6581, CP => CLK_I, Q => 
                           n_1378, QN => n4204);
   KEY_EXPAN0_reg_55_30_inst : FD1 port map( D => n6580, CP => CLK_I, Q => 
                           n_1379, QN => n4191);
   KEY_EXPAN0_reg_54_30_inst : FD1 port map( D => n6579, CP => CLK_I, Q => 
                           n_1380, QN => n4190);
   KEY_EXPAN0_reg_53_30_inst : FD1 port map( D => n6578, CP => CLK_I, Q => 
                           n_1381, QN => n4193);
   KEY_EXPAN0_reg_52_30_inst : FD1 port map( D => n6577, CP => CLK_I, Q => 
                           n_1382, QN => n4192);
   KEY_EXPAN0_reg_51_30_inst : FD1 port map( D => n6576, CP => CLK_I, Q => 
                           n_1383, QN => n4195);
   KEY_EXPAN0_reg_50_30_inst : FD1 port map( D => n6575, CP => CLK_I, Q => 
                           n_1384, QN => n4194);
   KEY_EXPAN0_reg_49_30_inst : FD1 port map( D => n6574, CP => CLK_I, Q => 
                           n_1385, QN => n4197);
   KEY_EXPAN0_reg_48_30_inst : FD1 port map( D => n6573, CP => CLK_I, Q => 
                           n_1386, QN => n4196);
   KEY_EXPAN0_reg_47_30_inst : FD1 port map( D => n6572, CP => CLK_I, Q => 
                           n_1387, QN => n4183);
   KEY_EXPAN0_reg_46_30_inst : FD1 port map( D => n6571, CP => CLK_I, Q => 
                           n_1388, QN => n4182);
   KEY_EXPAN0_reg_45_30_inst : FD1 port map( D => n6570, CP => CLK_I, Q => 
                           n_1389, QN => n4185);
   KEY_EXPAN0_reg_44_30_inst : FD1 port map( D => n6569, CP => CLK_I, Q => 
                           n_1390, QN => n4184);
   KEY_EXPAN0_reg_43_30_inst : FD1 port map( D => n6568, CP => CLK_I, Q => 
                           n_1391, QN => n4187);
   KEY_EXPAN0_reg_42_30_inst : FD1 port map( D => n6567, CP => CLK_I, Q => 
                           n_1392, QN => n4186);
   KEY_EXPAN0_reg_41_30_inst : FD1 port map( D => n6566, CP => CLK_I, Q => 
                           n_1393, QN => n4189);
   KEY_EXPAN0_reg_40_30_inst : FD1 port map( D => n6565, CP => CLK_I, Q => 
                           n_1394, QN => n4188);
   KEY_EXPAN0_reg_39_30_inst : FD1 port map( D => n6564, CP => CLK_I, Q => 
                           n_1395, QN => n4175);
   KEY_EXPAN0_reg_38_30_inst : FD1 port map( D => n6563, CP => CLK_I, Q => 
                           n_1396, QN => n4174);
   KEY_EXPAN0_reg_37_30_inst : FD1 port map( D => n6562, CP => CLK_I, Q => 
                           n_1397, QN => n4177);
   KEY_EXPAN0_reg_36_30_inst : FD1 port map( D => n6561, CP => CLK_I, Q => 
                           n_1398, QN => n4176);
   KEY_EXPAN0_reg_35_30_inst : FD1 port map( D => n6560, CP => CLK_I, Q => 
                           n_1399, QN => n4179);
   KEY_EXPAN0_reg_34_30_inst : FD1 port map( D => n6559, CP => CLK_I, Q => 
                           n_1400, QN => n4178);
   KEY_EXPAN0_reg_33_30_inst : FD1 port map( D => n6558, CP => CLK_I, Q => 
                           n_1401, QN => n4181);
   KEY_EXPAN0_reg_32_30_inst : FD1 port map( D => n6557, CP => CLK_I, Q => 
                           n_1402, QN => n4180);
   KEY_EXPAN0_reg_31_30_inst : FD1 port map( D => n6556, CP => CLK_I, Q => 
                           n_1403, QN => n4231);
   KEY_EXPAN0_reg_30_30_inst : FD1 port map( D => n6555, CP => CLK_I, Q => 
                           n_1404, QN => n4230);
   KEY_EXPAN0_reg_29_30_inst : FD1 port map( D => n6554, CP => CLK_I, Q => 
                           n_1405, QN => n4233);
   KEY_EXPAN0_reg_28_30_inst : FD1 port map( D => n6553, CP => CLK_I, Q => 
                           n_1406, QN => n4232);
   KEY_EXPAN0_reg_27_30_inst : FD1 port map( D => n6552, CP => CLK_I, Q => 
                           n_1407, QN => n4235);
   KEY_EXPAN0_reg_26_30_inst : FD1 port map( D => n6551, CP => CLK_I, Q => 
                           n_1408, QN => n4234);
   KEY_EXPAN0_reg_25_30_inst : FD1 port map( D => n6550, CP => CLK_I, Q => 
                           n_1409, QN => n4237);
   KEY_EXPAN0_reg_24_30_inst : FD1 port map( D => n6549, CP => CLK_I, Q => 
                           n_1410, QN => n4236);
   KEY_EXPAN0_reg_23_30_inst : FD1 port map( D => n6548, CP => CLK_I, Q => 
                           n_1411, QN => n4223);
   KEY_EXPAN0_reg_22_30_inst : FD1 port map( D => n6547, CP => CLK_I, Q => 
                           n_1412, QN => n4222);
   KEY_EXPAN0_reg_21_30_inst : FD1 port map( D => n6546, CP => CLK_I, Q => 
                           n_1413, QN => n4225);
   KEY_EXPAN0_reg_20_30_inst : FD1 port map( D => n6545, CP => CLK_I, Q => 
                           n_1414, QN => n4224);
   KEY_EXPAN0_reg_19_30_inst : FD1 port map( D => n6544, CP => CLK_I, Q => 
                           n_1415, QN => n4227);
   KEY_EXPAN0_reg_18_30_inst : FD1 port map( D => n6543, CP => CLK_I, Q => 
                           n_1416, QN => n4226);
   KEY_EXPAN0_reg_17_30_inst : FD1 port map( D => n6542, CP => CLK_I, Q => 
                           n_1417, QN => n4229);
   KEY_EXPAN0_reg_16_30_inst : FD1 port map( D => n6541, CP => CLK_I, Q => 
                           n_1418, QN => n4228);
   KEY_EXPAN0_reg_15_30_inst : FD1 port map( D => n6540, CP => CLK_I, Q => 
                           n_1419, QN => n4215);
   KEY_EXPAN0_reg_14_30_inst : FD1 port map( D => n6539, CP => CLK_I, Q => 
                           n_1420, QN => n4214);
   KEY_EXPAN0_reg_13_30_inst : FD1 port map( D => n6538, CP => CLK_I, Q => 
                           n_1421, QN => n4217);
   KEY_EXPAN0_reg_12_30_inst : FD1 port map( D => n6537, CP => CLK_I, Q => 
                           n_1422, QN => n4216);
   KEY_EXPAN0_reg_11_30_inst : FD1 port map( D => n6536, CP => CLK_I, Q => 
                           n_1423, QN => n4219);
   KEY_EXPAN0_reg_10_30_inst : FD1 port map( D => n6535, CP => CLK_I, Q => 
                           n_1424, QN => n4218);
   KEY_EXPAN0_reg_9_30_inst : FD1 port map( D => n6534, CP => CLK_I, Q => 
                           n_1425, QN => n4221);
   KEY_EXPAN0_reg_8_30_inst : FD1 port map( D => n6533, CP => CLK_I, Q => 
                           n_1426, QN => n4220);
   KEY_EXPAN0_reg_7_30_inst : FD1 port map( D => n6532, CP => CLK_I, Q => 
                           n_1427, QN => n4207);
   KEY_EXPAN0_reg_6_30_inst : FD1 port map( D => n6531, CP => CLK_I, Q => 
                           n_1428, QN => n4206);
   KEY_EXPAN0_reg_5_30_inst : FD1 port map( D => n6530, CP => CLK_I, Q => 
                           n_1429, QN => n4209);
   KEY_EXPAN0_reg_4_30_inst : FD1 port map( D => n6529, CP => CLK_I, Q => 
                           n_1430, QN => n4208);
   KEY_EXPAN0_reg_3_30_inst : FD1 port map( D => n6528, CP => CLK_I, Q => 
                           n_1431, QN => n4211);
   KEY_EXPAN0_reg_2_30_inst : FD1 port map( D => n6527, CP => CLK_I, Q => 
                           n_1432, QN => n4210);
   KEY_EXPAN0_reg_1_30_inst : FD1 port map( D => n6526, CP => CLK_I, Q => 
                           n_1433, QN => n4213);
   KEY_EXPAN0_reg_0_30_inst : FD1 port map( D => n6525, CP => CLK_I, Q => 
                           n_1434, QN => n4212);
   v_KEY_COL_OUT0_reg_30_inst : FD1 port map( D => n4590, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_30_port, QN => n1865);
   v_TEMP_VECTOR_reg_22_inst : FD1 port map( D => n6687, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_22_port, QN => n_1435);
   KEY_EXPAN0_reg_63_22_inst : FD1 port map( D => n6076, CP => CLK_I, Q => 
                           n_1436, QN => n4135);
   KEY_EXPAN0_reg_62_22_inst : FD1 port map( D => n6075, CP => CLK_I, Q => 
                           n_1437, QN => n4134);
   KEY_EXPAN0_reg_61_22_inst : FD1 port map( D => n6074, CP => CLK_I, Q => 
                           n_1438, QN => n4137);
   KEY_EXPAN0_reg_60_22_inst : FD1 port map( D => n6073, CP => CLK_I, Q => 
                           n_1439, QN => n4136);
   KEY_EXPAN0_reg_59_22_inst : FD1 port map( D => n6072, CP => CLK_I, Q => 
                           n_1440, QN => n4139);
   KEY_EXPAN0_reg_58_22_inst : FD1 port map( D => n6071, CP => CLK_I, Q => 
                           n_1441, QN => n4138);
   KEY_EXPAN0_reg_57_22_inst : FD1 port map( D => n6070, CP => CLK_I, Q => 
                           n_1442, QN => n4141);
   KEY_EXPAN0_reg_56_22_inst : FD1 port map( D => n6069, CP => CLK_I, Q => 
                           n_1443, QN => n4140);
   KEY_EXPAN0_reg_55_22_inst : FD1 port map( D => n6068, CP => CLK_I, Q => 
                           n_1444, QN => n4127);
   KEY_EXPAN0_reg_54_22_inst : FD1 port map( D => n6067, CP => CLK_I, Q => 
                           n_1445, QN => n4126);
   KEY_EXPAN0_reg_53_22_inst : FD1 port map( D => n6066, CP => CLK_I, Q => 
                           n_1446, QN => n4129);
   KEY_EXPAN0_reg_52_22_inst : FD1 port map( D => n6065, CP => CLK_I, Q => 
                           n_1447, QN => n4128);
   KEY_EXPAN0_reg_51_22_inst : FD1 port map( D => n6064, CP => CLK_I, Q => 
                           n_1448, QN => n4131);
   KEY_EXPAN0_reg_50_22_inst : FD1 port map( D => n6063, CP => CLK_I, Q => 
                           n_1449, QN => n4130);
   KEY_EXPAN0_reg_49_22_inst : FD1 port map( D => n6062, CP => CLK_I, Q => 
                           n_1450, QN => n4133);
   KEY_EXPAN0_reg_48_22_inst : FD1 port map( D => n6061, CP => CLK_I, Q => 
                           n_1451, QN => n4132);
   KEY_EXPAN0_reg_47_22_inst : FD1 port map( D => n6060, CP => CLK_I, Q => 
                           n_1452, QN => n4119);
   KEY_EXPAN0_reg_46_22_inst : FD1 port map( D => n6059, CP => CLK_I, Q => 
                           n_1453, QN => n4118);
   KEY_EXPAN0_reg_45_22_inst : FD1 port map( D => n6058, CP => CLK_I, Q => 
                           n_1454, QN => n4121);
   KEY_EXPAN0_reg_44_22_inst : FD1 port map( D => n6057, CP => CLK_I, Q => 
                           n_1455, QN => n4120);
   KEY_EXPAN0_reg_43_22_inst : FD1 port map( D => n6056, CP => CLK_I, Q => 
                           n_1456, QN => n4123);
   KEY_EXPAN0_reg_42_22_inst : FD1 port map( D => n6055, CP => CLK_I, Q => 
                           n_1457, QN => n4122);
   KEY_EXPAN0_reg_41_22_inst : FD1 port map( D => n6054, CP => CLK_I, Q => 
                           n_1458, QN => n4125);
   KEY_EXPAN0_reg_40_22_inst : FD1 port map( D => n6053, CP => CLK_I, Q => 
                           n_1459, QN => n4124);
   KEY_EXPAN0_reg_39_22_inst : FD1 port map( D => n6052, CP => CLK_I, Q => 
                           n_1460, QN => n4111);
   KEY_EXPAN0_reg_38_22_inst : FD1 port map( D => n6051, CP => CLK_I, Q => 
                           n_1461, QN => n4110);
   KEY_EXPAN0_reg_37_22_inst : FD1 port map( D => n6050, CP => CLK_I, Q => 
                           n_1462, QN => n4113);
   KEY_EXPAN0_reg_36_22_inst : FD1 port map( D => n6049, CP => CLK_I, Q => 
                           n_1463, QN => n4112);
   KEY_EXPAN0_reg_35_22_inst : FD1 port map( D => n6048, CP => CLK_I, Q => 
                           n_1464, QN => n4115);
   KEY_EXPAN0_reg_34_22_inst : FD1 port map( D => n6047, CP => CLK_I, Q => 
                           n_1465, QN => n4114);
   KEY_EXPAN0_reg_33_22_inst : FD1 port map( D => n6046, CP => CLK_I, Q => 
                           n_1466, QN => n4117);
   KEY_EXPAN0_reg_32_22_inst : FD1 port map( D => n6045, CP => CLK_I, Q => 
                           n_1467, QN => n4116);
   KEY_EXPAN0_reg_31_22_inst : FD1 port map( D => n6044, CP => CLK_I, Q => 
                           n_1468, QN => n4167);
   KEY_EXPAN0_reg_30_22_inst : FD1 port map( D => n6043, CP => CLK_I, Q => 
                           n_1469, QN => n4166);
   KEY_EXPAN0_reg_29_22_inst : FD1 port map( D => n6042, CP => CLK_I, Q => 
                           n_1470, QN => n4169);
   KEY_EXPAN0_reg_28_22_inst : FD1 port map( D => n6041, CP => CLK_I, Q => 
                           n_1471, QN => n4168);
   KEY_EXPAN0_reg_27_22_inst : FD1 port map( D => n6040, CP => CLK_I, Q => 
                           n_1472, QN => n4171);
   KEY_EXPAN0_reg_26_22_inst : FD1 port map( D => n6039, CP => CLK_I, Q => 
                           n_1473, QN => n4170);
   KEY_EXPAN0_reg_25_22_inst : FD1 port map( D => n6038, CP => CLK_I, Q => 
                           n_1474, QN => n4173);
   KEY_EXPAN0_reg_24_22_inst : FD1 port map( D => n6037, CP => CLK_I, Q => 
                           n_1475, QN => n4172);
   KEY_EXPAN0_reg_23_22_inst : FD1 port map( D => n6036, CP => CLK_I, Q => 
                           n_1476, QN => n4159);
   KEY_EXPAN0_reg_22_22_inst : FD1 port map( D => n6035, CP => CLK_I, Q => 
                           n_1477, QN => n4158);
   KEY_EXPAN0_reg_21_22_inst : FD1 port map( D => n6034, CP => CLK_I, Q => 
                           n_1478, QN => n4161);
   KEY_EXPAN0_reg_20_22_inst : FD1 port map( D => n6033, CP => CLK_I, Q => 
                           n_1479, QN => n4160);
   KEY_EXPAN0_reg_19_22_inst : FD1 port map( D => n6032, CP => CLK_I, Q => 
                           n_1480, QN => n4163);
   KEY_EXPAN0_reg_18_22_inst : FD1 port map( D => n6031, CP => CLK_I, Q => 
                           n_1481, QN => n4162);
   KEY_EXPAN0_reg_17_22_inst : FD1 port map( D => n6030, CP => CLK_I, Q => 
                           n_1482, QN => n4165);
   KEY_EXPAN0_reg_16_22_inst : FD1 port map( D => n6029, CP => CLK_I, Q => 
                           n_1483, QN => n4164);
   KEY_EXPAN0_reg_15_22_inst : FD1 port map( D => n6028, CP => CLK_I, Q => 
                           n_1484, QN => n4151);
   KEY_EXPAN0_reg_14_22_inst : FD1 port map( D => n6027, CP => CLK_I, Q => 
                           n_1485, QN => n4150);
   KEY_EXPAN0_reg_13_22_inst : FD1 port map( D => n6026, CP => CLK_I, Q => 
                           n_1486, QN => n4153);
   KEY_EXPAN0_reg_12_22_inst : FD1 port map( D => n6025, CP => CLK_I, Q => 
                           n_1487, QN => n4152);
   KEY_EXPAN0_reg_11_22_inst : FD1 port map( D => n6024, CP => CLK_I, Q => 
                           n_1488, QN => n4155);
   KEY_EXPAN0_reg_10_22_inst : FD1 port map( D => n6023, CP => CLK_I, Q => 
                           n_1489, QN => n4154);
   KEY_EXPAN0_reg_9_22_inst : FD1 port map( D => n6022, CP => CLK_I, Q => 
                           n_1490, QN => n4157);
   KEY_EXPAN0_reg_8_22_inst : FD1 port map( D => n6021, CP => CLK_I, Q => 
                           n_1491, QN => n4156);
   KEY_EXPAN0_reg_7_22_inst : FD1 port map( D => n6020, CP => CLK_I, Q => 
                           n_1492, QN => n4143);
   KEY_EXPAN0_reg_6_22_inst : FD1 port map( D => n6019, CP => CLK_I, Q => 
                           n_1493, QN => n4142);
   KEY_EXPAN0_reg_5_22_inst : FD1 port map( D => n6018, CP => CLK_I, Q => 
                           n_1494, QN => n4145);
   KEY_EXPAN0_reg_4_22_inst : FD1 port map( D => n6017, CP => CLK_I, Q => 
                           n_1495, QN => n4144);
   KEY_EXPAN0_reg_3_22_inst : FD1 port map( D => n6016, CP => CLK_I, Q => 
                           n_1496, QN => n4147);
   KEY_EXPAN0_reg_2_22_inst : FD1 port map( D => n6015, CP => CLK_I, Q => 
                           n_1497, QN => n4146);
   KEY_EXPAN0_reg_1_22_inst : FD1 port map( D => n6014, CP => CLK_I, Q => 
                           n_1498, QN => n4149);
   KEY_EXPAN0_reg_0_22_inst : FD1 port map( D => n6013, CP => CLK_I, Q => 
                           n_1499, QN => n4148);
   v_KEY_COL_OUT0_reg_22_inst : FD1 port map( D => n4589, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_22_port, QN => n1910);
   v_TEMP_VECTOR_reg_14_inst : FD1 port map( D => n6695, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_14_port, QN => n_1500);
   KEY_EXPAN0_reg_63_14_inst : FD1 port map( D => n5564, CP => CLK_I, Q => 
                           n_1501, QN => n4071);
   KEY_EXPAN0_reg_62_14_inst : FD1 port map( D => n5563, CP => CLK_I, Q => 
                           n_1502, QN => n4070);
   KEY_EXPAN0_reg_61_14_inst : FD1 port map( D => n5562, CP => CLK_I, Q => 
                           n_1503, QN => n4073);
   KEY_EXPAN0_reg_60_14_inst : FD1 port map( D => n5561, CP => CLK_I, Q => 
                           n_1504, QN => n4072);
   KEY_EXPAN0_reg_59_14_inst : FD1 port map( D => n5560, CP => CLK_I, Q => 
                           n_1505, QN => n4075);
   KEY_EXPAN0_reg_58_14_inst : FD1 port map( D => n5559, CP => CLK_I, Q => 
                           n_1506, QN => n4074);
   KEY_EXPAN0_reg_57_14_inst : FD1 port map( D => n5558, CP => CLK_I, Q => 
                           n_1507, QN => n4077);
   KEY_EXPAN0_reg_56_14_inst : FD1 port map( D => n5557, CP => CLK_I, Q => 
                           n_1508, QN => n4076);
   KEY_EXPAN0_reg_55_14_inst : FD1 port map( D => n5556, CP => CLK_I, Q => 
                           n_1509, QN => n4063);
   KEY_EXPAN0_reg_54_14_inst : FD1 port map( D => n5555, CP => CLK_I, Q => 
                           n_1510, QN => n4062);
   KEY_EXPAN0_reg_53_14_inst : FD1 port map( D => n5554, CP => CLK_I, Q => 
                           n_1511, QN => n4065);
   KEY_EXPAN0_reg_52_14_inst : FD1 port map( D => n5553, CP => CLK_I, Q => 
                           n_1512, QN => n4064);
   KEY_EXPAN0_reg_51_14_inst : FD1 port map( D => n5552, CP => CLK_I, Q => 
                           n_1513, QN => n4067);
   KEY_EXPAN0_reg_50_14_inst : FD1 port map( D => n5551, CP => CLK_I, Q => 
                           n_1514, QN => n4066);
   KEY_EXPAN0_reg_49_14_inst : FD1 port map( D => n5550, CP => CLK_I, Q => 
                           n_1515, QN => n4069);
   KEY_EXPAN0_reg_48_14_inst : FD1 port map( D => n5549, CP => CLK_I, Q => 
                           n_1516, QN => n4068);
   KEY_EXPAN0_reg_47_14_inst : FD1 port map( D => n5548, CP => CLK_I, Q => 
                           n_1517, QN => n4055);
   KEY_EXPAN0_reg_46_14_inst : FD1 port map( D => n5547, CP => CLK_I, Q => 
                           n_1518, QN => n4054);
   KEY_EXPAN0_reg_45_14_inst : FD1 port map( D => n5546, CP => CLK_I, Q => 
                           n_1519, QN => n4057);
   KEY_EXPAN0_reg_44_14_inst : FD1 port map( D => n5545, CP => CLK_I, Q => 
                           n_1520, QN => n4056);
   KEY_EXPAN0_reg_43_14_inst : FD1 port map( D => n5544, CP => CLK_I, Q => 
                           n_1521, QN => n4059);
   KEY_EXPAN0_reg_42_14_inst : FD1 port map( D => n5543, CP => CLK_I, Q => 
                           n_1522, QN => n4058);
   KEY_EXPAN0_reg_41_14_inst : FD1 port map( D => n5542, CP => CLK_I, Q => 
                           n_1523, QN => n4061);
   KEY_EXPAN0_reg_40_14_inst : FD1 port map( D => n5541, CP => CLK_I, Q => 
                           n_1524, QN => n4060);
   KEY_EXPAN0_reg_39_14_inst : FD1 port map( D => n5540, CP => CLK_I, Q => 
                           n_1525, QN => n4047);
   KEY_EXPAN0_reg_38_14_inst : FD1 port map( D => n5539, CP => CLK_I, Q => 
                           n_1526, QN => n4046);
   KEY_EXPAN0_reg_37_14_inst : FD1 port map( D => n5538, CP => CLK_I, Q => 
                           n_1527, QN => n4049);
   KEY_EXPAN0_reg_36_14_inst : FD1 port map( D => n5537, CP => CLK_I, Q => 
                           n_1528, QN => n4048);
   KEY_EXPAN0_reg_35_14_inst : FD1 port map( D => n5536, CP => CLK_I, Q => 
                           n_1529, QN => n4051);
   KEY_EXPAN0_reg_34_14_inst : FD1 port map( D => n5535, CP => CLK_I, Q => 
                           n_1530, QN => n4050);
   KEY_EXPAN0_reg_33_14_inst : FD1 port map( D => n5534, CP => CLK_I, Q => 
                           n_1531, QN => n4053);
   KEY_EXPAN0_reg_32_14_inst : FD1 port map( D => n5533, CP => CLK_I, Q => 
                           n_1532, QN => n4052);
   KEY_EXPAN0_reg_31_14_inst : FD1 port map( D => n5532, CP => CLK_I, Q => 
                           n_1533, QN => n4103);
   KEY_EXPAN0_reg_30_14_inst : FD1 port map( D => n5531, CP => CLK_I, Q => 
                           n_1534, QN => n4102);
   KEY_EXPAN0_reg_29_14_inst : FD1 port map( D => n5530, CP => CLK_I, Q => 
                           n_1535, QN => n4105);
   KEY_EXPAN0_reg_28_14_inst : FD1 port map( D => n5529, CP => CLK_I, Q => 
                           n_1536, QN => n4104);
   KEY_EXPAN0_reg_27_14_inst : FD1 port map( D => n5528, CP => CLK_I, Q => 
                           n_1537, QN => n4107);
   KEY_EXPAN0_reg_26_14_inst : FD1 port map( D => n5527, CP => CLK_I, Q => 
                           n_1538, QN => n4106);
   KEY_EXPAN0_reg_25_14_inst : FD1 port map( D => n5526, CP => CLK_I, Q => 
                           n_1539, QN => n4109);
   KEY_EXPAN0_reg_24_14_inst : FD1 port map( D => n5525, CP => CLK_I, Q => 
                           n_1540, QN => n4108);
   KEY_EXPAN0_reg_23_14_inst : FD1 port map( D => n5524, CP => CLK_I, Q => 
                           n_1541, QN => n4095);
   KEY_EXPAN0_reg_22_14_inst : FD1 port map( D => n5523, CP => CLK_I, Q => 
                           n_1542, QN => n4094);
   KEY_EXPAN0_reg_21_14_inst : FD1 port map( D => n5522, CP => CLK_I, Q => 
                           n_1543, QN => n4097);
   KEY_EXPAN0_reg_20_14_inst : FD1 port map( D => n5521, CP => CLK_I, Q => 
                           n_1544, QN => n4096);
   KEY_EXPAN0_reg_19_14_inst : FD1 port map( D => n5520, CP => CLK_I, Q => 
                           n_1545, QN => n4099);
   KEY_EXPAN0_reg_18_14_inst : FD1 port map( D => n5519, CP => CLK_I, Q => 
                           n_1546, QN => n4098);
   KEY_EXPAN0_reg_17_14_inst : FD1 port map( D => n5518, CP => CLK_I, Q => 
                           n_1547, QN => n4101);
   KEY_EXPAN0_reg_16_14_inst : FD1 port map( D => n5517, CP => CLK_I, Q => 
                           n_1548, QN => n4100);
   KEY_EXPAN0_reg_15_14_inst : FD1 port map( D => n5516, CP => CLK_I, Q => 
                           n_1549, QN => n4087);
   KEY_EXPAN0_reg_14_14_inst : FD1 port map( D => n5515, CP => CLK_I, Q => 
                           n_1550, QN => n4086);
   KEY_EXPAN0_reg_13_14_inst : FD1 port map( D => n5514, CP => CLK_I, Q => 
                           n_1551, QN => n4089);
   KEY_EXPAN0_reg_12_14_inst : FD1 port map( D => n5513, CP => CLK_I, Q => 
                           n_1552, QN => n4088);
   KEY_EXPAN0_reg_11_14_inst : FD1 port map( D => n5512, CP => CLK_I, Q => 
                           n_1553, QN => n4091);
   KEY_EXPAN0_reg_10_14_inst : FD1 port map( D => n5511, CP => CLK_I, Q => 
                           n_1554, QN => n4090);
   KEY_EXPAN0_reg_9_14_inst : FD1 port map( D => n5510, CP => CLK_I, Q => 
                           n_1555, QN => n4093);
   KEY_EXPAN0_reg_8_14_inst : FD1 port map( D => n5509, CP => CLK_I, Q => 
                           n_1556, QN => n4092);
   KEY_EXPAN0_reg_7_14_inst : FD1 port map( D => n5508, CP => CLK_I, Q => 
                           n_1557, QN => n4079);
   KEY_EXPAN0_reg_6_14_inst : FD1 port map( D => n5507, CP => CLK_I, Q => 
                           n_1558, QN => n4078);
   KEY_EXPAN0_reg_5_14_inst : FD1 port map( D => n5506, CP => CLK_I, Q => 
                           n_1559, QN => n4081);
   KEY_EXPAN0_reg_4_14_inst : FD1 port map( D => n5505, CP => CLK_I, Q => 
                           n_1560, QN => n4080);
   KEY_EXPAN0_reg_3_14_inst : FD1 port map( D => n5504, CP => CLK_I, Q => 
                           n_1561, QN => n4083);
   KEY_EXPAN0_reg_2_14_inst : FD1 port map( D => n5503, CP => CLK_I, Q => 
                           n_1562, QN => n4082);
   KEY_EXPAN0_reg_1_14_inst : FD1 port map( D => n5502, CP => CLK_I, Q => 
                           n_1563, QN => n4085);
   KEY_EXPAN0_reg_0_14_inst : FD1 port map( D => n5501, CP => CLK_I, Q => 
                           n_1564, QN => n4084);
   v_KEY_COL_OUT0_reg_14_inst : FD1 port map( D => n4588, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_14_port, QN => n1862);
   v_TEMP_VECTOR_reg_5_inst : FD1 port map( D => n6704, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_5_port, QN => n_1565);
   KEY_EXPAN0_reg_63_5_inst : FD1 port map( D => n4988, CP => CLK_I, Q => 
                           n_1566, QN => n4007);
   KEY_EXPAN0_reg_62_5_inst : FD1 port map( D => n4987, CP => CLK_I, Q => 
                           n_1567, QN => n4006);
   KEY_EXPAN0_reg_61_5_inst : FD1 port map( D => n4986, CP => CLK_I, Q => 
                           n_1568, QN => n4009);
   KEY_EXPAN0_reg_60_5_inst : FD1 port map( D => n4985, CP => CLK_I, Q => 
                           n_1569, QN => n4008);
   KEY_EXPAN0_reg_59_5_inst : FD1 port map( D => n4984, CP => CLK_I, Q => 
                           n_1570, QN => n4011);
   KEY_EXPAN0_reg_58_5_inst : FD1 port map( D => n4983, CP => CLK_I, Q => 
                           n_1571, QN => n4010);
   KEY_EXPAN0_reg_57_5_inst : FD1 port map( D => n4982, CP => CLK_I, Q => 
                           n_1572, QN => n4013);
   KEY_EXPAN0_reg_56_5_inst : FD1 port map( D => n4981, CP => CLK_I, Q => 
                           n_1573, QN => n4012);
   KEY_EXPAN0_reg_55_5_inst : FD1 port map( D => n4980, CP => CLK_I, Q => 
                           n_1574, QN => n3999);
   KEY_EXPAN0_reg_54_5_inst : FD1 port map( D => n4979, CP => CLK_I, Q => 
                           n_1575, QN => n3998);
   KEY_EXPAN0_reg_53_5_inst : FD1 port map( D => n4978, CP => CLK_I, Q => 
                           n_1576, QN => n4001);
   KEY_EXPAN0_reg_52_5_inst : FD1 port map( D => n4977, CP => CLK_I, Q => 
                           n_1577, QN => n4000);
   KEY_EXPAN0_reg_51_5_inst : FD1 port map( D => n4976, CP => CLK_I, Q => 
                           n_1578, QN => n4003);
   KEY_EXPAN0_reg_50_5_inst : FD1 port map( D => n4975, CP => CLK_I, Q => 
                           n_1579, QN => n4002);
   KEY_EXPAN0_reg_49_5_inst : FD1 port map( D => n4974, CP => CLK_I, Q => 
                           n_1580, QN => n4005);
   KEY_EXPAN0_reg_48_5_inst : FD1 port map( D => n4973, CP => CLK_I, Q => 
                           n_1581, QN => n4004);
   KEY_EXPAN0_reg_47_5_inst : FD1 port map( D => n4972, CP => CLK_I, Q => 
                           n_1582, QN => n3991);
   KEY_EXPAN0_reg_46_5_inst : FD1 port map( D => n4971, CP => CLK_I, Q => 
                           n_1583, QN => n3990);
   KEY_EXPAN0_reg_45_5_inst : FD1 port map( D => n4970, CP => CLK_I, Q => 
                           n_1584, QN => n3993);
   KEY_EXPAN0_reg_44_5_inst : FD1 port map( D => n4969, CP => CLK_I, Q => 
                           n_1585, QN => n3992);
   KEY_EXPAN0_reg_43_5_inst : FD1 port map( D => n4968, CP => CLK_I, Q => 
                           n_1586, QN => n3995);
   KEY_EXPAN0_reg_42_5_inst : FD1 port map( D => n4967, CP => CLK_I, Q => 
                           n_1587, QN => n3994);
   KEY_EXPAN0_reg_41_5_inst : FD1 port map( D => n4966, CP => CLK_I, Q => 
                           n_1588, QN => n3997);
   KEY_EXPAN0_reg_40_5_inst : FD1 port map( D => n4965, CP => CLK_I, Q => 
                           n_1589, QN => n3996);
   KEY_EXPAN0_reg_39_5_inst : FD1 port map( D => n4964, CP => CLK_I, Q => 
                           n_1590, QN => n3983);
   KEY_EXPAN0_reg_38_5_inst : FD1 port map( D => n4963, CP => CLK_I, Q => 
                           n_1591, QN => n3982);
   KEY_EXPAN0_reg_37_5_inst : FD1 port map( D => n4962, CP => CLK_I, Q => 
                           n_1592, QN => n3985);
   KEY_EXPAN0_reg_36_5_inst : FD1 port map( D => n4961, CP => CLK_I, Q => 
                           n_1593, QN => n3984);
   KEY_EXPAN0_reg_35_5_inst : FD1 port map( D => n4960, CP => CLK_I, Q => 
                           n_1594, QN => n3987);
   KEY_EXPAN0_reg_34_5_inst : FD1 port map( D => n4959, CP => CLK_I, Q => 
                           n_1595, QN => n3986);
   KEY_EXPAN0_reg_33_5_inst : FD1 port map( D => n4958, CP => CLK_I, Q => 
                           n_1596, QN => n3989);
   KEY_EXPAN0_reg_32_5_inst : FD1 port map( D => n4957, CP => CLK_I, Q => 
                           n_1597, QN => n3988);
   KEY_EXPAN0_reg_31_5_inst : FD1 port map( D => n4956, CP => CLK_I, Q => 
                           n_1598, QN => n4039);
   KEY_EXPAN0_reg_30_5_inst : FD1 port map( D => n4955, CP => CLK_I, Q => 
                           n_1599, QN => n4038);
   KEY_EXPAN0_reg_29_5_inst : FD1 port map( D => n4954, CP => CLK_I, Q => 
                           n_1600, QN => n4041);
   KEY_EXPAN0_reg_28_5_inst : FD1 port map( D => n4953, CP => CLK_I, Q => 
                           n_1601, QN => n4040);
   KEY_EXPAN0_reg_27_5_inst : FD1 port map( D => n4952, CP => CLK_I, Q => 
                           n_1602, QN => n4043);
   KEY_EXPAN0_reg_26_5_inst : FD1 port map( D => n4951, CP => CLK_I, Q => 
                           n_1603, QN => n4042);
   KEY_EXPAN0_reg_25_5_inst : FD1 port map( D => n4950, CP => CLK_I, Q => 
                           n_1604, QN => n4045);
   KEY_EXPAN0_reg_24_5_inst : FD1 port map( D => n4949, CP => CLK_I, Q => 
                           n_1605, QN => n4044);
   KEY_EXPAN0_reg_23_5_inst : FD1 port map( D => n4948, CP => CLK_I, Q => 
                           n_1606, QN => n4031);
   KEY_EXPAN0_reg_22_5_inst : FD1 port map( D => n4947, CP => CLK_I, Q => 
                           n_1607, QN => n4030);
   KEY_EXPAN0_reg_21_5_inst : FD1 port map( D => n4946, CP => CLK_I, Q => 
                           n_1608, QN => n4033);
   KEY_EXPAN0_reg_20_5_inst : FD1 port map( D => n4945, CP => CLK_I, Q => 
                           n_1609, QN => n4032);
   KEY_EXPAN0_reg_19_5_inst : FD1 port map( D => n4944, CP => CLK_I, Q => 
                           n_1610, QN => n4035);
   KEY_EXPAN0_reg_18_5_inst : FD1 port map( D => n4943, CP => CLK_I, Q => 
                           n_1611, QN => n4034);
   KEY_EXPAN0_reg_17_5_inst : FD1 port map( D => n4942, CP => CLK_I, Q => 
                           n_1612, QN => n4037);
   KEY_EXPAN0_reg_16_5_inst : FD1 port map( D => n4941, CP => CLK_I, Q => 
                           n_1613, QN => n4036);
   KEY_EXPAN0_reg_15_5_inst : FD1 port map( D => n4940, CP => CLK_I, Q => 
                           n_1614, QN => n4023);
   KEY_EXPAN0_reg_14_5_inst : FD1 port map( D => n4939, CP => CLK_I, Q => 
                           n_1615, QN => n4022);
   KEY_EXPAN0_reg_13_5_inst : FD1 port map( D => n4938, CP => CLK_I, Q => 
                           n_1616, QN => n4025);
   KEY_EXPAN0_reg_12_5_inst : FD1 port map( D => n4937, CP => CLK_I, Q => 
                           n_1617, QN => n4024);
   KEY_EXPAN0_reg_11_5_inst : FD1 port map( D => n4936, CP => CLK_I, Q => 
                           n_1618, QN => n4027);
   KEY_EXPAN0_reg_10_5_inst : FD1 port map( D => n4935, CP => CLK_I, Q => 
                           n_1619, QN => n4026);
   KEY_EXPAN0_reg_9_5_inst : FD1 port map( D => n4934, CP => CLK_I, Q => n_1620
                           , QN => n4029);
   KEY_EXPAN0_reg_8_5_inst : FD1 port map( D => n4933, CP => CLK_I, Q => n_1621
                           , QN => n4028);
   KEY_EXPAN0_reg_7_5_inst : FD1 port map( D => n4932, CP => CLK_I, Q => n_1622
                           , QN => n4015);
   KEY_EXPAN0_reg_6_5_inst : FD1 port map( D => n4931, CP => CLK_I, Q => n_1623
                           , QN => n4014);
   KEY_EXPAN0_reg_5_5_inst : FD1 port map( D => n4930, CP => CLK_I, Q => n_1624
                           , QN => n4017);
   KEY_EXPAN0_reg_4_5_inst : FD1 port map( D => n4929, CP => CLK_I, Q => n_1625
                           , QN => n4016);
   KEY_EXPAN0_reg_3_5_inst : FD1 port map( D => n4928, CP => CLK_I, Q => n_1626
                           , QN => n4019);
   KEY_EXPAN0_reg_2_5_inst : FD1 port map( D => n4927, CP => CLK_I, Q => n_1627
                           , QN => n4018);
   KEY_EXPAN0_reg_1_5_inst : FD1 port map( D => n4926, CP => CLK_I, Q => n_1628
                           , QN => n4021);
   KEY_EXPAN0_reg_0_5_inst : FD1 port map( D => n4925, CP => CLK_I, Q => n_1629
                           , QN => n4020);
   v_KEY_COL_OUT0_reg_5_inst : FD1 port map( D => n4587, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_5_port, QN => n1906);
   v_TEMP_VECTOR_reg_29_inst : FD1 port map( D => n6680, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_29_port, QN => n_1630);
   KEY_EXPAN0_reg_63_29_inst : FD1 port map( D => n6524, CP => CLK_I, Q => 
                           n_1631, QN => n3943);
   KEY_EXPAN0_reg_62_29_inst : FD1 port map( D => n6523, CP => CLK_I, Q => 
                           n_1632, QN => n3942);
   KEY_EXPAN0_reg_61_29_inst : FD1 port map( D => n6522, CP => CLK_I, Q => 
                           n_1633, QN => n3945);
   KEY_EXPAN0_reg_60_29_inst : FD1 port map( D => n6521, CP => CLK_I, Q => 
                           n_1634, QN => n3944);
   KEY_EXPAN0_reg_59_29_inst : FD1 port map( D => n6520, CP => CLK_I, Q => 
                           n_1635, QN => n3947);
   KEY_EXPAN0_reg_58_29_inst : FD1 port map( D => n6519, CP => CLK_I, Q => 
                           n_1636, QN => n3946);
   KEY_EXPAN0_reg_57_29_inst : FD1 port map( D => n6518, CP => CLK_I, Q => 
                           n_1637, QN => n3949);
   KEY_EXPAN0_reg_56_29_inst : FD1 port map( D => n6517, CP => CLK_I, Q => 
                           n_1638, QN => n3948);
   KEY_EXPAN0_reg_55_29_inst : FD1 port map( D => n6516, CP => CLK_I, Q => 
                           n_1639, QN => n3935);
   KEY_EXPAN0_reg_54_29_inst : FD1 port map( D => n6515, CP => CLK_I, Q => 
                           n_1640, QN => n3934);
   KEY_EXPAN0_reg_53_29_inst : FD1 port map( D => n6514, CP => CLK_I, Q => 
                           n_1641, QN => n3937);
   KEY_EXPAN0_reg_52_29_inst : FD1 port map( D => n6513, CP => CLK_I, Q => 
                           n_1642, QN => n3936);
   KEY_EXPAN0_reg_51_29_inst : FD1 port map( D => n6512, CP => CLK_I, Q => 
                           n_1643, QN => n3939);
   KEY_EXPAN0_reg_50_29_inst : FD1 port map( D => n6511, CP => CLK_I, Q => 
                           n_1644, QN => n3938);
   KEY_EXPAN0_reg_49_29_inst : FD1 port map( D => n6510, CP => CLK_I, Q => 
                           n_1645, QN => n3941);
   KEY_EXPAN0_reg_48_29_inst : FD1 port map( D => n6509, CP => CLK_I, Q => 
                           n_1646, QN => n3940);
   KEY_EXPAN0_reg_47_29_inst : FD1 port map( D => n6508, CP => CLK_I, Q => 
                           n_1647, QN => n3927);
   KEY_EXPAN0_reg_46_29_inst : FD1 port map( D => n6507, CP => CLK_I, Q => 
                           n_1648, QN => n3926);
   KEY_EXPAN0_reg_45_29_inst : FD1 port map( D => n6506, CP => CLK_I, Q => 
                           n_1649, QN => n3929);
   KEY_EXPAN0_reg_44_29_inst : FD1 port map( D => n6505, CP => CLK_I, Q => 
                           n_1650, QN => n3928);
   KEY_EXPAN0_reg_43_29_inst : FD1 port map( D => n6504, CP => CLK_I, Q => 
                           n_1651, QN => n3931);
   KEY_EXPAN0_reg_42_29_inst : FD1 port map( D => n6503, CP => CLK_I, Q => 
                           n_1652, QN => n3930);
   KEY_EXPAN0_reg_41_29_inst : FD1 port map( D => n6502, CP => CLK_I, Q => 
                           n_1653, QN => n3933);
   KEY_EXPAN0_reg_40_29_inst : FD1 port map( D => n6501, CP => CLK_I, Q => 
                           n_1654, QN => n3932);
   KEY_EXPAN0_reg_39_29_inst : FD1 port map( D => n6500, CP => CLK_I, Q => 
                           n_1655, QN => n3919);
   KEY_EXPAN0_reg_38_29_inst : FD1 port map( D => n6499, CP => CLK_I, Q => 
                           n_1656, QN => n3918);
   KEY_EXPAN0_reg_37_29_inst : FD1 port map( D => n6498, CP => CLK_I, Q => 
                           n_1657, QN => n3921);
   KEY_EXPAN0_reg_36_29_inst : FD1 port map( D => n6497, CP => CLK_I, Q => 
                           n_1658, QN => n3920);
   KEY_EXPAN0_reg_35_29_inst : FD1 port map( D => n6496, CP => CLK_I, Q => 
                           n_1659, QN => n3923);
   KEY_EXPAN0_reg_34_29_inst : FD1 port map( D => n6495, CP => CLK_I, Q => 
                           n_1660, QN => n3922);
   KEY_EXPAN0_reg_33_29_inst : FD1 port map( D => n6494, CP => CLK_I, Q => 
                           n_1661, QN => n3925);
   KEY_EXPAN0_reg_32_29_inst : FD1 port map( D => n6493, CP => CLK_I, Q => 
                           n_1662, QN => n3924);
   KEY_EXPAN0_reg_31_29_inst : FD1 port map( D => n6492, CP => CLK_I, Q => 
                           n_1663, QN => n3975);
   KEY_EXPAN0_reg_30_29_inst : FD1 port map( D => n6491, CP => CLK_I, Q => 
                           n_1664, QN => n3974);
   KEY_EXPAN0_reg_29_29_inst : FD1 port map( D => n6490, CP => CLK_I, Q => 
                           n_1665, QN => n3977);
   KEY_EXPAN0_reg_28_29_inst : FD1 port map( D => n6489, CP => CLK_I, Q => 
                           n_1666, QN => n3976);
   KEY_EXPAN0_reg_27_29_inst : FD1 port map( D => n6488, CP => CLK_I, Q => 
                           n_1667, QN => n3979);
   KEY_EXPAN0_reg_26_29_inst : FD1 port map( D => n6487, CP => CLK_I, Q => 
                           n_1668, QN => n3978);
   KEY_EXPAN0_reg_25_29_inst : FD1 port map( D => n6486, CP => CLK_I, Q => 
                           n_1669, QN => n3981);
   KEY_EXPAN0_reg_24_29_inst : FD1 port map( D => n6485, CP => CLK_I, Q => 
                           n_1670, QN => n3980);
   KEY_EXPAN0_reg_23_29_inst : FD1 port map( D => n6484, CP => CLK_I, Q => 
                           n_1671, QN => n3967);
   KEY_EXPAN0_reg_22_29_inst : FD1 port map( D => n6483, CP => CLK_I, Q => 
                           n_1672, QN => n3966);
   KEY_EXPAN0_reg_21_29_inst : FD1 port map( D => n6482, CP => CLK_I, Q => 
                           n_1673, QN => n3969);
   KEY_EXPAN0_reg_20_29_inst : FD1 port map( D => n6481, CP => CLK_I, Q => 
                           n_1674, QN => n3968);
   KEY_EXPAN0_reg_19_29_inst : FD1 port map( D => n6480, CP => CLK_I, Q => 
                           n_1675, QN => n3971);
   KEY_EXPAN0_reg_18_29_inst : FD1 port map( D => n6479, CP => CLK_I, Q => 
                           n_1676, QN => n3970);
   KEY_EXPAN0_reg_17_29_inst : FD1 port map( D => n6478, CP => CLK_I, Q => 
                           n_1677, QN => n3973);
   KEY_EXPAN0_reg_16_29_inst : FD1 port map( D => n6477, CP => CLK_I, Q => 
                           n_1678, QN => n3972);
   KEY_EXPAN0_reg_15_29_inst : FD1 port map( D => n6476, CP => CLK_I, Q => 
                           n_1679, QN => n3959);
   KEY_EXPAN0_reg_14_29_inst : FD1 port map( D => n6475, CP => CLK_I, Q => 
                           n_1680, QN => n3958);
   KEY_EXPAN0_reg_13_29_inst : FD1 port map( D => n6474, CP => CLK_I, Q => 
                           n_1681, QN => n3961);
   KEY_EXPAN0_reg_12_29_inst : FD1 port map( D => n6473, CP => CLK_I, Q => 
                           n_1682, QN => n3960);
   KEY_EXPAN0_reg_11_29_inst : FD1 port map( D => n6472, CP => CLK_I, Q => 
                           n_1683, QN => n3963);
   KEY_EXPAN0_reg_10_29_inst : FD1 port map( D => n6471, CP => CLK_I, Q => 
                           n_1684, QN => n3962);
   KEY_EXPAN0_reg_9_29_inst : FD1 port map( D => n6470, CP => CLK_I, Q => 
                           n_1685, QN => n3965);
   KEY_EXPAN0_reg_8_29_inst : FD1 port map( D => n6469, CP => CLK_I, Q => 
                           n_1686, QN => n3964);
   KEY_EXPAN0_reg_7_29_inst : FD1 port map( D => n6468, CP => CLK_I, Q => 
                           n_1687, QN => n3951);
   KEY_EXPAN0_reg_6_29_inst : FD1 port map( D => n6467, CP => CLK_I, Q => 
                           n_1688, QN => n3950);
   KEY_EXPAN0_reg_5_29_inst : FD1 port map( D => n6466, CP => CLK_I, Q => 
                           n_1689, QN => n3953);
   KEY_EXPAN0_reg_4_29_inst : FD1 port map( D => n6465, CP => CLK_I, Q => 
                           n_1690, QN => n3952);
   KEY_EXPAN0_reg_3_29_inst : FD1 port map( D => n6464, CP => CLK_I, Q => 
                           n_1691, QN => n3955);
   KEY_EXPAN0_reg_2_29_inst : FD1 port map( D => n6463, CP => CLK_I, Q => 
                           n_1692, QN => n3954);
   KEY_EXPAN0_reg_1_29_inst : FD1 port map( D => n6462, CP => CLK_I, Q => 
                           n_1693, QN => n3957);
   KEY_EXPAN0_reg_0_29_inst : FD1 port map( D => n6461, CP => CLK_I, Q => 
                           n_1694, QN => n3956);
   v_KEY_COL_OUT0_reg_29_inst : FD1 port map( D => n4586, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_29_port, QN => n1921);
   v_TEMP_VECTOR_reg_21_inst : FD1 port map( D => n6688, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_21_port, QN => n_1695);
   KEY_EXPAN0_reg_63_21_inst : FD1 port map( D => n6012, CP => CLK_I, Q => 
                           n_1696, QN => n3879);
   KEY_EXPAN0_reg_62_21_inst : FD1 port map( D => n6011, CP => CLK_I, Q => 
                           n_1697, QN => n3878);
   KEY_EXPAN0_reg_61_21_inst : FD1 port map( D => n6010, CP => CLK_I, Q => 
                           n_1698, QN => n3881);
   KEY_EXPAN0_reg_60_21_inst : FD1 port map( D => n6009, CP => CLK_I, Q => 
                           n_1699, QN => n3880);
   KEY_EXPAN0_reg_59_21_inst : FD1 port map( D => n6008, CP => CLK_I, Q => 
                           n_1700, QN => n3883);
   KEY_EXPAN0_reg_58_21_inst : FD1 port map( D => n6007, CP => CLK_I, Q => 
                           n_1701, QN => n3882);
   KEY_EXPAN0_reg_57_21_inst : FD1 port map( D => n6006, CP => CLK_I, Q => 
                           n_1702, QN => n3885);
   KEY_EXPAN0_reg_56_21_inst : FD1 port map( D => n6005, CP => CLK_I, Q => 
                           n_1703, QN => n3884);
   KEY_EXPAN0_reg_55_21_inst : FD1 port map( D => n6004, CP => CLK_I, Q => 
                           n_1704, QN => n3871);
   KEY_EXPAN0_reg_54_21_inst : FD1 port map( D => n6003, CP => CLK_I, Q => 
                           n_1705, QN => n3870);
   KEY_EXPAN0_reg_53_21_inst : FD1 port map( D => n6002, CP => CLK_I, Q => 
                           n_1706, QN => n3873);
   KEY_EXPAN0_reg_52_21_inst : FD1 port map( D => n6001, CP => CLK_I, Q => 
                           n_1707, QN => n3872);
   KEY_EXPAN0_reg_51_21_inst : FD1 port map( D => n6000, CP => CLK_I, Q => 
                           n_1708, QN => n3875);
   KEY_EXPAN0_reg_50_21_inst : FD1 port map( D => n5999, CP => CLK_I, Q => 
                           n_1709, QN => n3874);
   KEY_EXPAN0_reg_49_21_inst : FD1 port map( D => n5998, CP => CLK_I, Q => 
                           n_1710, QN => n3877);
   KEY_EXPAN0_reg_48_21_inst : FD1 port map( D => n5997, CP => CLK_I, Q => 
                           n_1711, QN => n3876);
   KEY_EXPAN0_reg_47_21_inst : FD1 port map( D => n5996, CP => CLK_I, Q => 
                           n_1712, QN => n3863);
   KEY_EXPAN0_reg_46_21_inst : FD1 port map( D => n5995, CP => CLK_I, Q => 
                           n_1713, QN => n3862);
   KEY_EXPAN0_reg_45_21_inst : FD1 port map( D => n5994, CP => CLK_I, Q => 
                           n_1714, QN => n3865);
   KEY_EXPAN0_reg_44_21_inst : FD1 port map( D => n5993, CP => CLK_I, Q => 
                           n_1715, QN => n3864);
   KEY_EXPAN0_reg_43_21_inst : FD1 port map( D => n5992, CP => CLK_I, Q => 
                           n_1716, QN => n3867);
   KEY_EXPAN0_reg_42_21_inst : FD1 port map( D => n5991, CP => CLK_I, Q => 
                           n_1717, QN => n3866);
   KEY_EXPAN0_reg_41_21_inst : FD1 port map( D => n5990, CP => CLK_I, Q => 
                           n_1718, QN => n3869);
   KEY_EXPAN0_reg_40_21_inst : FD1 port map( D => n5989, CP => CLK_I, Q => 
                           n_1719, QN => n3868);
   KEY_EXPAN0_reg_39_21_inst : FD1 port map( D => n5988, CP => CLK_I, Q => 
                           n_1720, QN => n3855);
   KEY_EXPAN0_reg_38_21_inst : FD1 port map( D => n5987, CP => CLK_I, Q => 
                           n_1721, QN => n3854);
   KEY_EXPAN0_reg_37_21_inst : FD1 port map( D => n5986, CP => CLK_I, Q => 
                           n_1722, QN => n3857);
   KEY_EXPAN0_reg_36_21_inst : FD1 port map( D => n5985, CP => CLK_I, Q => 
                           n_1723, QN => n3856);
   KEY_EXPAN0_reg_35_21_inst : FD1 port map( D => n5984, CP => CLK_I, Q => 
                           n_1724, QN => n3859);
   KEY_EXPAN0_reg_34_21_inst : FD1 port map( D => n5983, CP => CLK_I, Q => 
                           n_1725, QN => n3858);
   KEY_EXPAN0_reg_33_21_inst : FD1 port map( D => n5982, CP => CLK_I, Q => 
                           n_1726, QN => n3861);
   KEY_EXPAN0_reg_32_21_inst : FD1 port map( D => n5981, CP => CLK_I, Q => 
                           n_1727, QN => n3860);
   KEY_EXPAN0_reg_31_21_inst : FD1 port map( D => n5980, CP => CLK_I, Q => 
                           n_1728, QN => n3911);
   KEY_EXPAN0_reg_30_21_inst : FD1 port map( D => n5979, CP => CLK_I, Q => 
                           n_1729, QN => n3910);
   KEY_EXPAN0_reg_29_21_inst : FD1 port map( D => n5978, CP => CLK_I, Q => 
                           n_1730, QN => n3913);
   KEY_EXPAN0_reg_28_21_inst : FD1 port map( D => n5977, CP => CLK_I, Q => 
                           n_1731, QN => n3912);
   KEY_EXPAN0_reg_27_21_inst : FD1 port map( D => n5976, CP => CLK_I, Q => 
                           n_1732, QN => n3915);
   KEY_EXPAN0_reg_26_21_inst : FD1 port map( D => n5975, CP => CLK_I, Q => 
                           n_1733, QN => n3914);
   KEY_EXPAN0_reg_25_21_inst : FD1 port map( D => n5974, CP => CLK_I, Q => 
                           n_1734, QN => n3917);
   KEY_EXPAN0_reg_24_21_inst : FD1 port map( D => n5973, CP => CLK_I, Q => 
                           n_1735, QN => n3916);
   KEY_EXPAN0_reg_23_21_inst : FD1 port map( D => n5972, CP => CLK_I, Q => 
                           n_1736, QN => n3903);
   KEY_EXPAN0_reg_22_21_inst : FD1 port map( D => n5971, CP => CLK_I, Q => 
                           n_1737, QN => n3902);
   KEY_EXPAN0_reg_21_21_inst : FD1 port map( D => n5970, CP => CLK_I, Q => 
                           n_1738, QN => n3905);
   KEY_EXPAN0_reg_20_21_inst : FD1 port map( D => n5969, CP => CLK_I, Q => 
                           n_1739, QN => n3904);
   KEY_EXPAN0_reg_19_21_inst : FD1 port map( D => n5968, CP => CLK_I, Q => 
                           n_1740, QN => n3907);
   KEY_EXPAN0_reg_18_21_inst : FD1 port map( D => n5967, CP => CLK_I, Q => 
                           n_1741, QN => n3906);
   KEY_EXPAN0_reg_17_21_inst : FD1 port map( D => n5966, CP => CLK_I, Q => 
                           n_1742, QN => n3909);
   KEY_EXPAN0_reg_16_21_inst : FD1 port map( D => n5965, CP => CLK_I, Q => 
                           n_1743, QN => n3908);
   KEY_EXPAN0_reg_15_21_inst : FD1 port map( D => n5964, CP => CLK_I, Q => 
                           n_1744, QN => n3895);
   KEY_EXPAN0_reg_14_21_inst : FD1 port map( D => n5963, CP => CLK_I, Q => 
                           n_1745, QN => n3894);
   KEY_EXPAN0_reg_13_21_inst : FD1 port map( D => n5962, CP => CLK_I, Q => 
                           n_1746, QN => n3897);
   KEY_EXPAN0_reg_12_21_inst : FD1 port map( D => n5961, CP => CLK_I, Q => 
                           n_1747, QN => n3896);
   KEY_EXPAN0_reg_11_21_inst : FD1 port map( D => n5960, CP => CLK_I, Q => 
                           n_1748, QN => n3899);
   KEY_EXPAN0_reg_10_21_inst : FD1 port map( D => n5959, CP => CLK_I, Q => 
                           n_1749, QN => n3898);
   KEY_EXPAN0_reg_9_21_inst : FD1 port map( D => n5958, CP => CLK_I, Q => 
                           n_1750, QN => n3901);
   KEY_EXPAN0_reg_8_21_inst : FD1 port map( D => n5957, CP => CLK_I, Q => 
                           n_1751, QN => n3900);
   KEY_EXPAN0_reg_7_21_inst : FD1 port map( D => n5956, CP => CLK_I, Q => 
                           n_1752, QN => n3887);
   KEY_EXPAN0_reg_6_21_inst : FD1 port map( D => n5955, CP => CLK_I, Q => 
                           n_1753, QN => n3886);
   KEY_EXPAN0_reg_5_21_inst : FD1 port map( D => n5954, CP => CLK_I, Q => 
                           n_1754, QN => n3889);
   KEY_EXPAN0_reg_4_21_inst : FD1 port map( D => n5953, CP => CLK_I, Q => 
                           n_1755, QN => n3888);
   KEY_EXPAN0_reg_3_21_inst : FD1 port map( D => n5952, CP => CLK_I, Q => 
                           n_1756, QN => n3891);
   KEY_EXPAN0_reg_2_21_inst : FD1 port map( D => n5951, CP => CLK_I, Q => 
                           n_1757, QN => n3890);
   KEY_EXPAN0_reg_1_21_inst : FD1 port map( D => n5950, CP => CLK_I, Q => 
                           n_1758, QN => n3893);
   KEY_EXPAN0_reg_0_21_inst : FD1 port map( D => n5949, CP => CLK_I, Q => 
                           n_1759, QN => n3892);
   v_KEY_COL_OUT0_reg_21_inst : FD1 port map( D => n4585, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_21_port, QN => n1931);
   v_TEMP_VECTOR_reg_13_inst : FD1 port map( D => n6696, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_13_port, QN => n_1760);
   KEY_EXPAN0_reg_63_13_inst : FD1 port map( D => n5500, CP => CLK_I, Q => 
                           n_1761, QN => n3815);
   KEY_EXPAN0_reg_62_13_inst : FD1 port map( D => n5499, CP => CLK_I, Q => 
                           n_1762, QN => n3814);
   KEY_EXPAN0_reg_61_13_inst : FD1 port map( D => n5498, CP => CLK_I, Q => 
                           n_1763, QN => n3817);
   KEY_EXPAN0_reg_60_13_inst : FD1 port map( D => n5497, CP => CLK_I, Q => 
                           n_1764, QN => n3816);
   KEY_EXPAN0_reg_59_13_inst : FD1 port map( D => n5496, CP => CLK_I, Q => 
                           n_1765, QN => n3819);
   KEY_EXPAN0_reg_58_13_inst : FD1 port map( D => n5495, CP => CLK_I, Q => 
                           n_1766, QN => n3818);
   KEY_EXPAN0_reg_57_13_inst : FD1 port map( D => n5494, CP => CLK_I, Q => 
                           n_1767, QN => n3821);
   KEY_EXPAN0_reg_56_13_inst : FD1 port map( D => n5493, CP => CLK_I, Q => 
                           n_1768, QN => n3820);
   KEY_EXPAN0_reg_55_13_inst : FD1 port map( D => n5492, CP => CLK_I, Q => 
                           n_1769, QN => n3807);
   KEY_EXPAN0_reg_54_13_inst : FD1 port map( D => n5491, CP => CLK_I, Q => 
                           n_1770, QN => n3806);
   KEY_EXPAN0_reg_53_13_inst : FD1 port map( D => n5490, CP => CLK_I, Q => 
                           n_1771, QN => n3809);
   KEY_EXPAN0_reg_52_13_inst : FD1 port map( D => n5489, CP => CLK_I, Q => 
                           n_1772, QN => n3808);
   KEY_EXPAN0_reg_51_13_inst : FD1 port map( D => n5488, CP => CLK_I, Q => 
                           n_1773, QN => n3811);
   KEY_EXPAN0_reg_50_13_inst : FD1 port map( D => n5487, CP => CLK_I, Q => 
                           n_1774, QN => n3810);
   KEY_EXPAN0_reg_49_13_inst : FD1 port map( D => n5486, CP => CLK_I, Q => 
                           n_1775, QN => n3813);
   KEY_EXPAN0_reg_48_13_inst : FD1 port map( D => n5485, CP => CLK_I, Q => 
                           n_1776, QN => n3812);
   KEY_EXPAN0_reg_47_13_inst : FD1 port map( D => n5484, CP => CLK_I, Q => 
                           n_1777, QN => n3799);
   KEY_EXPAN0_reg_46_13_inst : FD1 port map( D => n5483, CP => CLK_I, Q => 
                           n_1778, QN => n3798);
   KEY_EXPAN0_reg_45_13_inst : FD1 port map( D => n5482, CP => CLK_I, Q => 
                           n_1779, QN => n3801);
   KEY_EXPAN0_reg_44_13_inst : FD1 port map( D => n5481, CP => CLK_I, Q => 
                           n_1780, QN => n3800);
   KEY_EXPAN0_reg_43_13_inst : FD1 port map( D => n5480, CP => CLK_I, Q => 
                           n_1781, QN => n3803);
   KEY_EXPAN0_reg_42_13_inst : FD1 port map( D => n5479, CP => CLK_I, Q => 
                           n_1782, QN => n3802);
   KEY_EXPAN0_reg_41_13_inst : FD1 port map( D => n5478, CP => CLK_I, Q => 
                           n_1783, QN => n3805);
   KEY_EXPAN0_reg_40_13_inst : FD1 port map( D => n5477, CP => CLK_I, Q => 
                           n_1784, QN => n3804);
   KEY_EXPAN0_reg_39_13_inst : FD1 port map( D => n5476, CP => CLK_I, Q => 
                           n_1785, QN => n3791);
   KEY_EXPAN0_reg_38_13_inst : FD1 port map( D => n5475, CP => CLK_I, Q => 
                           n_1786, QN => n3790);
   KEY_EXPAN0_reg_37_13_inst : FD1 port map( D => n5474, CP => CLK_I, Q => 
                           n_1787, QN => n3793);
   KEY_EXPAN0_reg_36_13_inst : FD1 port map( D => n5473, CP => CLK_I, Q => 
                           n_1788, QN => n3792);
   KEY_EXPAN0_reg_35_13_inst : FD1 port map( D => n5472, CP => CLK_I, Q => 
                           n_1789, QN => n3795);
   KEY_EXPAN0_reg_34_13_inst : FD1 port map( D => n5471, CP => CLK_I, Q => 
                           n_1790, QN => n3794);
   KEY_EXPAN0_reg_33_13_inst : FD1 port map( D => n5470, CP => CLK_I, Q => 
                           n_1791, QN => n3797);
   KEY_EXPAN0_reg_32_13_inst : FD1 port map( D => n5469, CP => CLK_I, Q => 
                           n_1792, QN => n3796);
   KEY_EXPAN0_reg_31_13_inst : FD1 port map( D => n5468, CP => CLK_I, Q => 
                           n_1793, QN => n3847);
   KEY_EXPAN0_reg_30_13_inst : FD1 port map( D => n5467, CP => CLK_I, Q => 
                           n_1794, QN => n3846);
   KEY_EXPAN0_reg_29_13_inst : FD1 port map( D => n5466, CP => CLK_I, Q => 
                           n_1795, QN => n3849);
   KEY_EXPAN0_reg_28_13_inst : FD1 port map( D => n5465, CP => CLK_I, Q => 
                           n_1796, QN => n3848);
   KEY_EXPAN0_reg_27_13_inst : FD1 port map( D => n5464, CP => CLK_I, Q => 
                           n_1797, QN => n3851);
   KEY_EXPAN0_reg_26_13_inst : FD1 port map( D => n5463, CP => CLK_I, Q => 
                           n_1798, QN => n3850);
   KEY_EXPAN0_reg_25_13_inst : FD1 port map( D => n5462, CP => CLK_I, Q => 
                           n_1799, QN => n3853);
   KEY_EXPAN0_reg_24_13_inst : FD1 port map( D => n5461, CP => CLK_I, Q => 
                           n_1800, QN => n3852);
   KEY_EXPAN0_reg_23_13_inst : FD1 port map( D => n5460, CP => CLK_I, Q => 
                           n_1801, QN => n3839);
   KEY_EXPAN0_reg_22_13_inst : FD1 port map( D => n5459, CP => CLK_I, Q => 
                           n_1802, QN => n3838);
   KEY_EXPAN0_reg_21_13_inst : FD1 port map( D => n5458, CP => CLK_I, Q => 
                           n_1803, QN => n3841);
   KEY_EXPAN0_reg_20_13_inst : FD1 port map( D => n5457, CP => CLK_I, Q => 
                           n_1804, QN => n3840);
   KEY_EXPAN0_reg_19_13_inst : FD1 port map( D => n5456, CP => CLK_I, Q => 
                           n_1805, QN => n3843);
   KEY_EXPAN0_reg_18_13_inst : FD1 port map( D => n5455, CP => CLK_I, Q => 
                           n_1806, QN => n3842);
   KEY_EXPAN0_reg_17_13_inst : FD1 port map( D => n5454, CP => CLK_I, Q => 
                           n_1807, QN => n3845);
   KEY_EXPAN0_reg_16_13_inst : FD1 port map( D => n5453, CP => CLK_I, Q => 
                           n_1808, QN => n3844);
   KEY_EXPAN0_reg_15_13_inst : FD1 port map( D => n5452, CP => CLK_I, Q => 
                           n_1809, QN => n3831);
   KEY_EXPAN0_reg_14_13_inst : FD1 port map( D => n5451, CP => CLK_I, Q => 
                           n_1810, QN => n3830);
   KEY_EXPAN0_reg_13_13_inst : FD1 port map( D => n5450, CP => CLK_I, Q => 
                           n_1811, QN => n3833);
   KEY_EXPAN0_reg_12_13_inst : FD1 port map( D => n5449, CP => CLK_I, Q => 
                           n_1812, QN => n3832);
   KEY_EXPAN0_reg_11_13_inst : FD1 port map( D => n5448, CP => CLK_I, Q => 
                           n_1813, QN => n3835);
   KEY_EXPAN0_reg_10_13_inst : FD1 port map( D => n5447, CP => CLK_I, Q => 
                           n_1814, QN => n3834);
   KEY_EXPAN0_reg_9_13_inst : FD1 port map( D => n5446, CP => CLK_I, Q => 
                           n_1815, QN => n3837);
   KEY_EXPAN0_reg_8_13_inst : FD1 port map( D => n5445, CP => CLK_I, Q => 
                           n_1816, QN => n3836);
   KEY_EXPAN0_reg_7_13_inst : FD1 port map( D => n5444, CP => CLK_I, Q => 
                           n_1817, QN => n3823);
   KEY_EXPAN0_reg_6_13_inst : FD1 port map( D => n5443, CP => CLK_I, Q => 
                           n_1818, QN => n3822);
   KEY_EXPAN0_reg_5_13_inst : FD1 port map( D => n5442, CP => CLK_I, Q => 
                           n_1819, QN => n3825);
   KEY_EXPAN0_reg_4_13_inst : FD1 port map( D => n5441, CP => CLK_I, Q => 
                           n_1820, QN => n3824);
   KEY_EXPAN0_reg_3_13_inst : FD1 port map( D => n5440, CP => CLK_I, Q => 
                           n_1821, QN => n3827);
   KEY_EXPAN0_reg_2_13_inst : FD1 port map( D => n5439, CP => CLK_I, Q => 
                           n_1822, QN => n3826);
   KEY_EXPAN0_reg_1_13_inst : FD1 port map( D => n5438, CP => CLK_I, Q => 
                           n_1823, QN => n3829);
   KEY_EXPAN0_reg_0_13_inst : FD1 port map( D => n5437, CP => CLK_I, Q => 
                           n_1824, QN => n3828);
   v_KEY_COL_OUT0_reg_13_inst : FD1 port map( D => n4584, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_13_port, QN => n1905);
   v_TEMP_VECTOR_reg_4_inst : FD1 port map( D => n6705, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_4_port, QN => n_1825);
   KEY_EXPAN0_reg_63_4_inst : FD1 port map( D => n4924, CP => CLK_I, Q => 
                           n_1826, QN => n3751);
   KEY_EXPAN0_reg_62_4_inst : FD1 port map( D => n4923, CP => CLK_I, Q => 
                           n_1827, QN => n3750);
   KEY_EXPAN0_reg_61_4_inst : FD1 port map( D => n4922, CP => CLK_I, Q => 
                           n_1828, QN => n3753);
   KEY_EXPAN0_reg_60_4_inst : FD1 port map( D => n4921, CP => CLK_I, Q => 
                           n_1829, QN => n3752);
   KEY_EXPAN0_reg_59_4_inst : FD1 port map( D => n4920, CP => CLK_I, Q => 
                           n_1830, QN => n3755);
   KEY_EXPAN0_reg_58_4_inst : FD1 port map( D => n4919, CP => CLK_I, Q => 
                           n_1831, QN => n3754);
   KEY_EXPAN0_reg_57_4_inst : FD1 port map( D => n4918, CP => CLK_I, Q => 
                           n_1832, QN => n3757);
   KEY_EXPAN0_reg_56_4_inst : FD1 port map( D => n4917, CP => CLK_I, Q => 
                           n_1833, QN => n3756);
   KEY_EXPAN0_reg_55_4_inst : FD1 port map( D => n4916, CP => CLK_I, Q => 
                           n_1834, QN => n3743);
   KEY_EXPAN0_reg_54_4_inst : FD1 port map( D => n4915, CP => CLK_I, Q => 
                           n_1835, QN => n3742);
   KEY_EXPAN0_reg_53_4_inst : FD1 port map( D => n4914, CP => CLK_I, Q => 
                           n_1836, QN => n3745);
   KEY_EXPAN0_reg_52_4_inst : FD1 port map( D => n4913, CP => CLK_I, Q => 
                           n_1837, QN => n3744);
   KEY_EXPAN0_reg_51_4_inst : FD1 port map( D => n4912, CP => CLK_I, Q => 
                           n_1838, QN => n3747);
   KEY_EXPAN0_reg_50_4_inst : FD1 port map( D => n4911, CP => CLK_I, Q => 
                           n_1839, QN => n3746);
   KEY_EXPAN0_reg_49_4_inst : FD1 port map( D => n4910, CP => CLK_I, Q => 
                           n_1840, QN => n3749);
   KEY_EXPAN0_reg_48_4_inst : FD1 port map( D => n4909, CP => CLK_I, Q => 
                           n_1841, QN => n3748);
   KEY_EXPAN0_reg_47_4_inst : FD1 port map( D => n4908, CP => CLK_I, Q => 
                           n_1842, QN => n3735);
   KEY_EXPAN0_reg_46_4_inst : FD1 port map( D => n4907, CP => CLK_I, Q => 
                           n_1843, QN => n3734);
   KEY_EXPAN0_reg_45_4_inst : FD1 port map( D => n4906, CP => CLK_I, Q => 
                           n_1844, QN => n3737);
   KEY_EXPAN0_reg_44_4_inst : FD1 port map( D => n4905, CP => CLK_I, Q => 
                           n_1845, QN => n3736);
   KEY_EXPAN0_reg_43_4_inst : FD1 port map( D => n4904, CP => CLK_I, Q => 
                           n_1846, QN => n3739);
   KEY_EXPAN0_reg_42_4_inst : FD1 port map( D => n4903, CP => CLK_I, Q => 
                           n_1847, QN => n3738);
   KEY_EXPAN0_reg_41_4_inst : FD1 port map( D => n4902, CP => CLK_I, Q => 
                           n_1848, QN => n3741);
   KEY_EXPAN0_reg_40_4_inst : FD1 port map( D => n4901, CP => CLK_I, Q => 
                           n_1849, QN => n3740);
   KEY_EXPAN0_reg_39_4_inst : FD1 port map( D => n4900, CP => CLK_I, Q => 
                           n_1850, QN => n3727);
   KEY_EXPAN0_reg_38_4_inst : FD1 port map( D => n4899, CP => CLK_I, Q => 
                           n_1851, QN => n3726);
   KEY_EXPAN0_reg_37_4_inst : FD1 port map( D => n4898, CP => CLK_I, Q => 
                           n_1852, QN => n3729);
   KEY_EXPAN0_reg_36_4_inst : FD1 port map( D => n4897, CP => CLK_I, Q => 
                           n_1853, QN => n3728);
   KEY_EXPAN0_reg_35_4_inst : FD1 port map( D => n4896, CP => CLK_I, Q => 
                           n_1854, QN => n3731);
   KEY_EXPAN0_reg_34_4_inst : FD1 port map( D => n4895, CP => CLK_I, Q => 
                           n_1855, QN => n3730);
   KEY_EXPAN0_reg_33_4_inst : FD1 port map( D => n4894, CP => CLK_I, Q => 
                           n_1856, QN => n3733);
   KEY_EXPAN0_reg_32_4_inst : FD1 port map( D => n4893, CP => CLK_I, Q => 
                           n_1857, QN => n3732);
   KEY_EXPAN0_reg_31_4_inst : FD1 port map( D => n4892, CP => CLK_I, Q => 
                           n_1858, QN => n3783);
   KEY_EXPAN0_reg_30_4_inst : FD1 port map( D => n4891, CP => CLK_I, Q => 
                           n_1859, QN => n3782);
   KEY_EXPAN0_reg_29_4_inst : FD1 port map( D => n4890, CP => CLK_I, Q => 
                           n_1860, QN => n3785);
   KEY_EXPAN0_reg_28_4_inst : FD1 port map( D => n4889, CP => CLK_I, Q => 
                           n_1861, QN => n3784);
   KEY_EXPAN0_reg_27_4_inst : FD1 port map( D => n4888, CP => CLK_I, Q => 
                           n_1862, QN => n3787);
   KEY_EXPAN0_reg_26_4_inst : FD1 port map( D => n4887, CP => CLK_I, Q => 
                           n_1863, QN => n3786);
   KEY_EXPAN0_reg_25_4_inst : FD1 port map( D => n4886, CP => CLK_I, Q => 
                           n_1864, QN => n3789);
   KEY_EXPAN0_reg_24_4_inst : FD1 port map( D => n4885, CP => CLK_I, Q => 
                           n_1865, QN => n3788);
   KEY_EXPAN0_reg_23_4_inst : FD1 port map( D => n4884, CP => CLK_I, Q => 
                           n_1866, QN => n3775);
   KEY_EXPAN0_reg_22_4_inst : FD1 port map( D => n4883, CP => CLK_I, Q => 
                           n_1867, QN => n3774);
   KEY_EXPAN0_reg_21_4_inst : FD1 port map( D => n4882, CP => CLK_I, Q => 
                           n_1868, QN => n3777);
   KEY_EXPAN0_reg_20_4_inst : FD1 port map( D => n4881, CP => CLK_I, Q => 
                           n_1869, QN => n3776);
   KEY_EXPAN0_reg_19_4_inst : FD1 port map( D => n4880, CP => CLK_I, Q => 
                           n_1870, QN => n3779);
   KEY_EXPAN0_reg_18_4_inst : FD1 port map( D => n4879, CP => CLK_I, Q => 
                           n_1871, QN => n3778);
   KEY_EXPAN0_reg_17_4_inst : FD1 port map( D => n4878, CP => CLK_I, Q => 
                           n_1872, QN => n3781);
   KEY_EXPAN0_reg_16_4_inst : FD1 port map( D => n4877, CP => CLK_I, Q => 
                           n_1873, QN => n3780);
   KEY_EXPAN0_reg_15_4_inst : FD1 port map( D => n4876, CP => CLK_I, Q => 
                           n_1874, QN => n3767);
   KEY_EXPAN0_reg_14_4_inst : FD1 port map( D => n4875, CP => CLK_I, Q => 
                           n_1875, QN => n3766);
   KEY_EXPAN0_reg_13_4_inst : FD1 port map( D => n4874, CP => CLK_I, Q => 
                           n_1876, QN => n3769);
   KEY_EXPAN0_reg_12_4_inst : FD1 port map( D => n4873, CP => CLK_I, Q => 
                           n_1877, QN => n3768);
   KEY_EXPAN0_reg_11_4_inst : FD1 port map( D => n4872, CP => CLK_I, Q => 
                           n_1878, QN => n3771);
   KEY_EXPAN0_reg_10_4_inst : FD1 port map( D => n4871, CP => CLK_I, Q => 
                           n_1879, QN => n3770);
   KEY_EXPAN0_reg_9_4_inst : FD1 port map( D => n4870, CP => CLK_I, Q => n_1880
                           , QN => n3773);
   KEY_EXPAN0_reg_8_4_inst : FD1 port map( D => n4869, CP => CLK_I, Q => n_1881
                           , QN => n3772);
   KEY_EXPAN0_reg_7_4_inst : FD1 port map( D => n4868, CP => CLK_I, Q => n_1882
                           , QN => n3759);
   KEY_EXPAN0_reg_6_4_inst : FD1 port map( D => n4867, CP => CLK_I, Q => n_1883
                           , QN => n3758);
   KEY_EXPAN0_reg_5_4_inst : FD1 port map( D => n4866, CP => CLK_I, Q => n_1884
                           , QN => n3761);
   KEY_EXPAN0_reg_4_4_inst : FD1 port map( D => n4865, CP => CLK_I, Q => n_1885
                           , QN => n3760);
   KEY_EXPAN0_reg_3_4_inst : FD1 port map( D => n4864, CP => CLK_I, Q => n_1886
                           , QN => n3763);
   KEY_EXPAN0_reg_2_4_inst : FD1 port map( D => n4863, CP => CLK_I, Q => n_1887
                           , QN => n3762);
   KEY_EXPAN0_reg_1_4_inst : FD1 port map( D => n4862, CP => CLK_I, Q => n_1888
                           , QN => n3765);
   KEY_EXPAN0_reg_0_4_inst : FD1 port map( D => n4861, CP => CLK_I, Q => n_1889
                           , QN => n3764);
   v_KEY_COL_OUT0_reg_4_inst : FD1 port map( D => n4583, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_4_port, QN => n2023);
   v_TEMP_VECTOR_reg_28_inst : FD1 port map( D => n6681, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_28_port, QN => n_1890);
   KEY_EXPAN0_reg_63_28_inst : FD1 port map( D => n6460, CP => CLK_I, Q => 
                           n_1891, QN => n3687);
   KEY_EXPAN0_reg_62_28_inst : FD1 port map( D => n6459, CP => CLK_I, Q => 
                           n_1892, QN => n3686);
   KEY_EXPAN0_reg_61_28_inst : FD1 port map( D => n6458, CP => CLK_I, Q => 
                           n_1893, QN => n3689);
   KEY_EXPAN0_reg_60_28_inst : FD1 port map( D => n6457, CP => CLK_I, Q => 
                           n_1894, QN => n3688);
   KEY_EXPAN0_reg_59_28_inst : FD1 port map( D => n6456, CP => CLK_I, Q => 
                           n_1895, QN => n3691);
   KEY_EXPAN0_reg_58_28_inst : FD1 port map( D => n6455, CP => CLK_I, Q => 
                           n_1896, QN => n3690);
   KEY_EXPAN0_reg_57_28_inst : FD1 port map( D => n6454, CP => CLK_I, Q => 
                           n_1897, QN => n3693);
   KEY_EXPAN0_reg_56_28_inst : FD1 port map( D => n6453, CP => CLK_I, Q => 
                           n_1898, QN => n3692);
   KEY_EXPAN0_reg_55_28_inst : FD1 port map( D => n6452, CP => CLK_I, Q => 
                           n_1899, QN => n3679);
   KEY_EXPAN0_reg_54_28_inst : FD1 port map( D => n6451, CP => CLK_I, Q => 
                           n_1900, QN => n3678);
   KEY_EXPAN0_reg_53_28_inst : FD1 port map( D => n6450, CP => CLK_I, Q => 
                           n_1901, QN => n3681);
   KEY_EXPAN0_reg_52_28_inst : FD1 port map( D => n6449, CP => CLK_I, Q => 
                           n_1902, QN => n3680);
   KEY_EXPAN0_reg_51_28_inst : FD1 port map( D => n6448, CP => CLK_I, Q => 
                           n_1903, QN => n3683);
   KEY_EXPAN0_reg_50_28_inst : FD1 port map( D => n6447, CP => CLK_I, Q => 
                           n_1904, QN => n3682);
   KEY_EXPAN0_reg_49_28_inst : FD1 port map( D => n6446, CP => CLK_I, Q => 
                           n_1905, QN => n3685);
   KEY_EXPAN0_reg_48_28_inst : FD1 port map( D => n6445, CP => CLK_I, Q => 
                           n_1906, QN => n3684);
   KEY_EXPAN0_reg_47_28_inst : FD1 port map( D => n6444, CP => CLK_I, Q => 
                           n_1907, QN => n3671);
   KEY_EXPAN0_reg_46_28_inst : FD1 port map( D => n6443, CP => CLK_I, Q => 
                           n_1908, QN => n3670);
   KEY_EXPAN0_reg_45_28_inst : FD1 port map( D => n6442, CP => CLK_I, Q => 
                           n_1909, QN => n3673);
   KEY_EXPAN0_reg_44_28_inst : FD1 port map( D => n6441, CP => CLK_I, Q => 
                           n_1910, QN => n3672);
   KEY_EXPAN0_reg_43_28_inst : FD1 port map( D => n6440, CP => CLK_I, Q => 
                           n_1911, QN => n3675);
   KEY_EXPAN0_reg_42_28_inst : FD1 port map( D => n6439, CP => CLK_I, Q => 
                           n_1912, QN => n3674);
   KEY_EXPAN0_reg_41_28_inst : FD1 port map( D => n6438, CP => CLK_I, Q => 
                           n_1913, QN => n3677);
   KEY_EXPAN0_reg_40_28_inst : FD1 port map( D => n6437, CP => CLK_I, Q => 
                           n_1914, QN => n3676);
   KEY_EXPAN0_reg_39_28_inst : FD1 port map( D => n6436, CP => CLK_I, Q => 
                           n_1915, QN => n3663);
   KEY_EXPAN0_reg_38_28_inst : FD1 port map( D => n6435, CP => CLK_I, Q => 
                           n_1916, QN => n3662);
   KEY_EXPAN0_reg_37_28_inst : FD1 port map( D => n6434, CP => CLK_I, Q => 
                           n_1917, QN => n3665);
   KEY_EXPAN0_reg_36_28_inst : FD1 port map( D => n6433, CP => CLK_I, Q => 
                           n_1918, QN => n3664);
   KEY_EXPAN0_reg_35_28_inst : FD1 port map( D => n6432, CP => CLK_I, Q => 
                           n_1919, QN => n3667);
   KEY_EXPAN0_reg_34_28_inst : FD1 port map( D => n6431, CP => CLK_I, Q => 
                           n_1920, QN => n3666);
   KEY_EXPAN0_reg_33_28_inst : FD1 port map( D => n6430, CP => CLK_I, Q => 
                           n_1921, QN => n3669);
   KEY_EXPAN0_reg_32_28_inst : FD1 port map( D => n6429, CP => CLK_I, Q => 
                           n_1922, QN => n3668);
   KEY_EXPAN0_reg_31_28_inst : FD1 port map( D => n6428, CP => CLK_I, Q => 
                           n_1923, QN => n3719);
   KEY_EXPAN0_reg_30_28_inst : FD1 port map( D => n6427, CP => CLK_I, Q => 
                           n_1924, QN => n3718);
   KEY_EXPAN0_reg_29_28_inst : FD1 port map( D => n6426, CP => CLK_I, Q => 
                           n_1925, QN => n3721);
   KEY_EXPAN0_reg_28_28_inst : FD1 port map( D => n6425, CP => CLK_I, Q => 
                           n_1926, QN => n3720);
   KEY_EXPAN0_reg_27_28_inst : FD1 port map( D => n6424, CP => CLK_I, Q => 
                           n_1927, QN => n3723);
   KEY_EXPAN0_reg_26_28_inst : FD1 port map( D => n6423, CP => CLK_I, Q => 
                           n_1928, QN => n3722);
   KEY_EXPAN0_reg_25_28_inst : FD1 port map( D => n6422, CP => CLK_I, Q => 
                           n_1929, QN => n3725);
   KEY_EXPAN0_reg_24_28_inst : FD1 port map( D => n6421, CP => CLK_I, Q => 
                           n_1930, QN => n3724);
   KEY_EXPAN0_reg_23_28_inst : FD1 port map( D => n6420, CP => CLK_I, Q => 
                           n_1931, QN => n3711);
   KEY_EXPAN0_reg_22_28_inst : FD1 port map( D => n6419, CP => CLK_I, Q => 
                           n_1932, QN => n3710);
   KEY_EXPAN0_reg_21_28_inst : FD1 port map( D => n6418, CP => CLK_I, Q => 
                           n_1933, QN => n3713);
   KEY_EXPAN0_reg_20_28_inst : FD1 port map( D => n6417, CP => CLK_I, Q => 
                           n_1934, QN => n3712);
   KEY_EXPAN0_reg_19_28_inst : FD1 port map( D => n6416, CP => CLK_I, Q => 
                           n_1935, QN => n3715);
   KEY_EXPAN0_reg_18_28_inst : FD1 port map( D => n6415, CP => CLK_I, Q => 
                           n_1936, QN => n3714);
   KEY_EXPAN0_reg_17_28_inst : FD1 port map( D => n6414, CP => CLK_I, Q => 
                           n_1937, QN => n3717);
   KEY_EXPAN0_reg_16_28_inst : FD1 port map( D => n6413, CP => CLK_I, Q => 
                           n_1938, QN => n3716);
   KEY_EXPAN0_reg_15_28_inst : FD1 port map( D => n6412, CP => CLK_I, Q => 
                           n_1939, QN => n3703);
   KEY_EXPAN0_reg_14_28_inst : FD1 port map( D => n6411, CP => CLK_I, Q => 
                           n_1940, QN => n3702);
   KEY_EXPAN0_reg_13_28_inst : FD1 port map( D => n6410, CP => CLK_I, Q => 
                           n_1941, QN => n3705);
   KEY_EXPAN0_reg_12_28_inst : FD1 port map( D => n6409, CP => CLK_I, Q => 
                           n_1942, QN => n3704);
   KEY_EXPAN0_reg_11_28_inst : FD1 port map( D => n6408, CP => CLK_I, Q => 
                           n_1943, QN => n3707);
   KEY_EXPAN0_reg_10_28_inst : FD1 port map( D => n6407, CP => CLK_I, Q => 
                           n_1944, QN => n3706);
   KEY_EXPAN0_reg_9_28_inst : FD1 port map( D => n6406, CP => CLK_I, Q => 
                           n_1945, QN => n3709);
   KEY_EXPAN0_reg_8_28_inst : FD1 port map( D => n6405, CP => CLK_I, Q => 
                           n_1946, QN => n3708);
   KEY_EXPAN0_reg_7_28_inst : FD1 port map( D => n6404, CP => CLK_I, Q => 
                           n_1947, QN => n3695);
   KEY_EXPAN0_reg_6_28_inst : FD1 port map( D => n6403, CP => CLK_I, Q => 
                           n_1948, QN => n3694);
   KEY_EXPAN0_reg_5_28_inst : FD1 port map( D => n6402, CP => CLK_I, Q => 
                           n_1949, QN => n3697);
   KEY_EXPAN0_reg_4_28_inst : FD1 port map( D => n6401, CP => CLK_I, Q => 
                           n_1950, QN => n3696);
   KEY_EXPAN0_reg_3_28_inst : FD1 port map( D => n6400, CP => CLK_I, Q => 
                           n_1951, QN => n3699);
   KEY_EXPAN0_reg_2_28_inst : FD1 port map( D => n6399, CP => CLK_I, Q => 
                           n_1952, QN => n3698);
   KEY_EXPAN0_reg_1_28_inst : FD1 port map( D => n6398, CP => CLK_I, Q => 
                           n_1953, QN => n3701);
   KEY_EXPAN0_reg_0_28_inst : FD1 port map( D => n6397, CP => CLK_I, Q => 
                           n_1954, QN => n3700);
   v_KEY_COL_OUT0_reg_28_inst : FD1 port map( D => n4582, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_28_port, QN => n1967);
   v_TEMP_VECTOR_reg_20_inst : FD1 port map( D => n6689, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_20_port, QN => n_1955);
   KEY_EXPAN0_reg_63_20_inst : FD1 port map( D => n5948, CP => CLK_I, Q => 
                           n_1956, QN => n3623);
   KEY_EXPAN0_reg_62_20_inst : FD1 port map( D => n5947, CP => CLK_I, Q => 
                           n_1957, QN => n3622);
   KEY_EXPAN0_reg_61_20_inst : FD1 port map( D => n5946, CP => CLK_I, Q => 
                           n_1958, QN => n3625);
   KEY_EXPAN0_reg_60_20_inst : FD1 port map( D => n5945, CP => CLK_I, Q => 
                           n_1959, QN => n3624);
   KEY_EXPAN0_reg_59_20_inst : FD1 port map( D => n5944, CP => CLK_I, Q => 
                           n_1960, QN => n3627);
   KEY_EXPAN0_reg_58_20_inst : FD1 port map( D => n5943, CP => CLK_I, Q => 
                           n_1961, QN => n3626);
   KEY_EXPAN0_reg_57_20_inst : FD1 port map( D => n5942, CP => CLK_I, Q => 
                           n_1962, QN => n3629);
   KEY_EXPAN0_reg_56_20_inst : FD1 port map( D => n5941, CP => CLK_I, Q => 
                           n_1963, QN => n3628);
   KEY_EXPAN0_reg_55_20_inst : FD1 port map( D => n5940, CP => CLK_I, Q => 
                           n_1964, QN => n3615);
   KEY_EXPAN0_reg_54_20_inst : FD1 port map( D => n5939, CP => CLK_I, Q => 
                           n_1965, QN => n3614);
   KEY_EXPAN0_reg_53_20_inst : FD1 port map( D => n5938, CP => CLK_I, Q => 
                           n_1966, QN => n3617);
   KEY_EXPAN0_reg_52_20_inst : FD1 port map( D => n5937, CP => CLK_I, Q => 
                           n_1967, QN => n3616);
   KEY_EXPAN0_reg_51_20_inst : FD1 port map( D => n5936, CP => CLK_I, Q => 
                           n_1968, QN => n3619);
   KEY_EXPAN0_reg_50_20_inst : FD1 port map( D => n5935, CP => CLK_I, Q => 
                           n_1969, QN => n3618);
   KEY_EXPAN0_reg_49_20_inst : FD1 port map( D => n5934, CP => CLK_I, Q => 
                           n_1970, QN => n3621);
   KEY_EXPAN0_reg_48_20_inst : FD1 port map( D => n5933, CP => CLK_I, Q => 
                           n_1971, QN => n3620);
   KEY_EXPAN0_reg_47_20_inst : FD1 port map( D => n5932, CP => CLK_I, Q => 
                           n_1972, QN => n3607);
   KEY_EXPAN0_reg_46_20_inst : FD1 port map( D => n5931, CP => CLK_I, Q => 
                           n_1973, QN => n3606);
   KEY_EXPAN0_reg_45_20_inst : FD1 port map( D => n5930, CP => CLK_I, Q => 
                           n_1974, QN => n3609);
   KEY_EXPAN0_reg_44_20_inst : FD1 port map( D => n5929, CP => CLK_I, Q => 
                           n_1975, QN => n3608);
   KEY_EXPAN0_reg_43_20_inst : FD1 port map( D => n5928, CP => CLK_I, Q => 
                           n_1976, QN => n3611);
   KEY_EXPAN0_reg_42_20_inst : FD1 port map( D => n5927, CP => CLK_I, Q => 
                           n_1977, QN => n3610);
   KEY_EXPAN0_reg_41_20_inst : FD1 port map( D => n5926, CP => CLK_I, Q => 
                           n_1978, QN => n3613);
   KEY_EXPAN0_reg_40_20_inst : FD1 port map( D => n5925, CP => CLK_I, Q => 
                           n_1979, QN => n3612);
   KEY_EXPAN0_reg_39_20_inst : FD1 port map( D => n5924, CP => CLK_I, Q => 
                           n_1980, QN => n3599);
   KEY_EXPAN0_reg_38_20_inst : FD1 port map( D => n5923, CP => CLK_I, Q => 
                           n_1981, QN => n3598);
   KEY_EXPAN0_reg_37_20_inst : FD1 port map( D => n5922, CP => CLK_I, Q => 
                           n_1982, QN => n3601);
   KEY_EXPAN0_reg_36_20_inst : FD1 port map( D => n5921, CP => CLK_I, Q => 
                           n_1983, QN => n3600);
   KEY_EXPAN0_reg_35_20_inst : FD1 port map( D => n5920, CP => CLK_I, Q => 
                           n_1984, QN => n3603);
   KEY_EXPAN0_reg_34_20_inst : FD1 port map( D => n5919, CP => CLK_I, Q => 
                           n_1985, QN => n3602);
   KEY_EXPAN0_reg_33_20_inst : FD1 port map( D => n5918, CP => CLK_I, Q => 
                           n_1986, QN => n3605);
   KEY_EXPAN0_reg_32_20_inst : FD1 port map( D => n5917, CP => CLK_I, Q => 
                           n_1987, QN => n3604);
   KEY_EXPAN0_reg_31_20_inst : FD1 port map( D => n5916, CP => CLK_I, Q => 
                           n_1988, QN => n3655);
   KEY_EXPAN0_reg_30_20_inst : FD1 port map( D => n5915, CP => CLK_I, Q => 
                           n_1989, QN => n3654);
   KEY_EXPAN0_reg_29_20_inst : FD1 port map( D => n5914, CP => CLK_I, Q => 
                           n_1990, QN => n3657);
   KEY_EXPAN0_reg_28_20_inst : FD1 port map( D => n5913, CP => CLK_I, Q => 
                           n_1991, QN => n3656);
   KEY_EXPAN0_reg_27_20_inst : FD1 port map( D => n5912, CP => CLK_I, Q => 
                           n_1992, QN => n3659);
   KEY_EXPAN0_reg_26_20_inst : FD1 port map( D => n5911, CP => CLK_I, Q => 
                           n_1993, QN => n3658);
   KEY_EXPAN0_reg_25_20_inst : FD1 port map( D => n5910, CP => CLK_I, Q => 
                           n_1994, QN => n3661);
   KEY_EXPAN0_reg_24_20_inst : FD1 port map( D => n5909, CP => CLK_I, Q => 
                           n_1995, QN => n3660);
   KEY_EXPAN0_reg_23_20_inst : FD1 port map( D => n5908, CP => CLK_I, Q => 
                           n_1996, QN => n3647);
   KEY_EXPAN0_reg_22_20_inst : FD1 port map( D => n5907, CP => CLK_I, Q => 
                           n_1997, QN => n3646);
   KEY_EXPAN0_reg_21_20_inst : FD1 port map( D => n5906, CP => CLK_I, Q => 
                           n_1998, QN => n3649);
   KEY_EXPAN0_reg_20_20_inst : FD1 port map( D => n5905, CP => CLK_I, Q => 
                           n_1999, QN => n3648);
   KEY_EXPAN0_reg_19_20_inst : FD1 port map( D => n5904, CP => CLK_I, Q => 
                           n_2000, QN => n3651);
   KEY_EXPAN0_reg_18_20_inst : FD1 port map( D => n5903, CP => CLK_I, Q => 
                           n_2001, QN => n3650);
   KEY_EXPAN0_reg_17_20_inst : FD1 port map( D => n5902, CP => CLK_I, Q => 
                           n_2002, QN => n3653);
   KEY_EXPAN0_reg_16_20_inst : FD1 port map( D => n5901, CP => CLK_I, Q => 
                           n_2003, QN => n3652);
   KEY_EXPAN0_reg_15_20_inst : FD1 port map( D => n5900, CP => CLK_I, Q => 
                           n_2004, QN => n3639);
   KEY_EXPAN0_reg_14_20_inst : FD1 port map( D => n5899, CP => CLK_I, Q => 
                           n_2005, QN => n3638);
   KEY_EXPAN0_reg_13_20_inst : FD1 port map( D => n5898, CP => CLK_I, Q => 
                           n_2006, QN => n3641);
   KEY_EXPAN0_reg_12_20_inst : FD1 port map( D => n5897, CP => CLK_I, Q => 
                           n_2007, QN => n3640);
   KEY_EXPAN0_reg_11_20_inst : FD1 port map( D => n5896, CP => CLK_I, Q => 
                           n_2008, QN => n3643);
   KEY_EXPAN0_reg_10_20_inst : FD1 port map( D => n5895, CP => CLK_I, Q => 
                           n_2009, QN => n3642);
   KEY_EXPAN0_reg_9_20_inst : FD1 port map( D => n5894, CP => CLK_I, Q => 
                           n_2010, QN => n3645);
   KEY_EXPAN0_reg_8_20_inst : FD1 port map( D => n5893, CP => CLK_I, Q => 
                           n_2011, QN => n3644);
   KEY_EXPAN0_reg_7_20_inst : FD1 port map( D => n5892, CP => CLK_I, Q => 
                           n_2012, QN => n3631);
   KEY_EXPAN0_reg_6_20_inst : FD1 port map( D => n5891, CP => CLK_I, Q => 
                           n_2013, QN => n3630);
   KEY_EXPAN0_reg_5_20_inst : FD1 port map( D => n5890, CP => CLK_I, Q => 
                           n_2014, QN => n3633);
   KEY_EXPAN0_reg_4_20_inst : FD1 port map( D => n5889, CP => CLK_I, Q => 
                           n_2015, QN => n3632);
   KEY_EXPAN0_reg_3_20_inst : FD1 port map( D => n5888, CP => CLK_I, Q => 
                           n_2016, QN => n3635);
   KEY_EXPAN0_reg_2_20_inst : FD1 port map( D => n5887, CP => CLK_I, Q => 
                           n_2017, QN => n3634);
   KEY_EXPAN0_reg_1_20_inst : FD1 port map( D => n5886, CP => CLK_I, Q => 
                           n_2018, QN => n3637);
   KEY_EXPAN0_reg_0_20_inst : FD1 port map( D => n5885, CP => CLK_I, Q => 
                           n_2019, QN => n3636);
   v_KEY_COL_OUT0_reg_20_inst : FD1 port map( D => n4581, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_20_port, QN => n1984);
   v_TEMP_VECTOR_reg_12_inst : FD1 port map( D => n6697, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_12_port, QN => n_2020);
   KEY_EXPAN0_reg_63_12_inst : FD1 port map( D => n5436, CP => CLK_I, Q => 
                           n_2021, QN => n3559);
   KEY_EXPAN0_reg_62_12_inst : FD1 port map( D => n5435, CP => CLK_I, Q => 
                           n_2022, QN => n3558);
   KEY_EXPAN0_reg_61_12_inst : FD1 port map( D => n5434, CP => CLK_I, Q => 
                           n_2023, QN => n3561);
   KEY_EXPAN0_reg_60_12_inst : FD1 port map( D => n5433, CP => CLK_I, Q => 
                           n_2024, QN => n3560);
   KEY_EXPAN0_reg_59_12_inst : FD1 port map( D => n5432, CP => CLK_I, Q => 
                           n_2025, QN => n3563);
   KEY_EXPAN0_reg_58_12_inst : FD1 port map( D => n5431, CP => CLK_I, Q => 
                           n_2026, QN => n3562);
   KEY_EXPAN0_reg_57_12_inst : FD1 port map( D => n5430, CP => CLK_I, Q => 
                           n_2027, QN => n3565);
   KEY_EXPAN0_reg_56_12_inst : FD1 port map( D => n5429, CP => CLK_I, Q => 
                           n_2028, QN => n3564);
   KEY_EXPAN0_reg_55_12_inst : FD1 port map( D => n5428, CP => CLK_I, Q => 
                           n_2029, QN => n3551);
   KEY_EXPAN0_reg_54_12_inst : FD1 port map( D => n5427, CP => CLK_I, Q => 
                           n_2030, QN => n3550);
   KEY_EXPAN0_reg_53_12_inst : FD1 port map( D => n5426, CP => CLK_I, Q => 
                           n_2031, QN => n3553);
   KEY_EXPAN0_reg_52_12_inst : FD1 port map( D => n5425, CP => CLK_I, Q => 
                           n_2032, QN => n3552);
   KEY_EXPAN0_reg_51_12_inst : FD1 port map( D => n5424, CP => CLK_I, Q => 
                           n_2033, QN => n3555);
   KEY_EXPAN0_reg_50_12_inst : FD1 port map( D => n5423, CP => CLK_I, Q => 
                           n_2034, QN => n3554);
   KEY_EXPAN0_reg_49_12_inst : FD1 port map( D => n5422, CP => CLK_I, Q => 
                           n_2035, QN => n3557);
   KEY_EXPAN0_reg_48_12_inst : FD1 port map( D => n5421, CP => CLK_I, Q => 
                           n_2036, QN => n3556);
   KEY_EXPAN0_reg_47_12_inst : FD1 port map( D => n5420, CP => CLK_I, Q => 
                           n_2037, QN => n3543);
   KEY_EXPAN0_reg_46_12_inst : FD1 port map( D => n5419, CP => CLK_I, Q => 
                           n_2038, QN => n3542);
   KEY_EXPAN0_reg_45_12_inst : FD1 port map( D => n5418, CP => CLK_I, Q => 
                           n_2039, QN => n3545);
   KEY_EXPAN0_reg_44_12_inst : FD1 port map( D => n5417, CP => CLK_I, Q => 
                           n_2040, QN => n3544);
   KEY_EXPAN0_reg_43_12_inst : FD1 port map( D => n5416, CP => CLK_I, Q => 
                           n_2041, QN => n3547);
   KEY_EXPAN0_reg_42_12_inst : FD1 port map( D => n5415, CP => CLK_I, Q => 
                           n_2042, QN => n3546);
   KEY_EXPAN0_reg_41_12_inst : FD1 port map( D => n5414, CP => CLK_I, Q => 
                           n_2043, QN => n3549);
   KEY_EXPAN0_reg_40_12_inst : FD1 port map( D => n5413, CP => CLK_I, Q => 
                           n_2044, QN => n3548);
   KEY_EXPAN0_reg_39_12_inst : FD1 port map( D => n5412, CP => CLK_I, Q => 
                           n_2045, QN => n3535);
   KEY_EXPAN0_reg_38_12_inst : FD1 port map( D => n5411, CP => CLK_I, Q => 
                           n_2046, QN => n3534);
   KEY_EXPAN0_reg_37_12_inst : FD1 port map( D => n5410, CP => CLK_I, Q => 
                           n_2047, QN => n3537);
   KEY_EXPAN0_reg_36_12_inst : FD1 port map( D => n5409, CP => CLK_I, Q => 
                           n_2048, QN => n3536);
   KEY_EXPAN0_reg_35_12_inst : FD1 port map( D => n5408, CP => CLK_I, Q => 
                           n_2049, QN => n3539);
   KEY_EXPAN0_reg_34_12_inst : FD1 port map( D => n5407, CP => CLK_I, Q => 
                           n_2050, QN => n3538);
   KEY_EXPAN0_reg_33_12_inst : FD1 port map( D => n5406, CP => CLK_I, Q => 
                           n_2051, QN => n3541);
   KEY_EXPAN0_reg_32_12_inst : FD1 port map( D => n5405, CP => CLK_I, Q => 
                           n_2052, QN => n3540);
   KEY_EXPAN0_reg_31_12_inst : FD1 port map( D => n5404, CP => CLK_I, Q => 
                           n_2053, QN => n3591);
   KEY_EXPAN0_reg_30_12_inst : FD1 port map( D => n5403, CP => CLK_I, Q => 
                           n_2054, QN => n3590);
   KEY_EXPAN0_reg_29_12_inst : FD1 port map( D => n5402, CP => CLK_I, Q => 
                           n_2055, QN => n3593);
   KEY_EXPAN0_reg_28_12_inst : FD1 port map( D => n5401, CP => CLK_I, Q => 
                           n_2056, QN => n3592);
   KEY_EXPAN0_reg_27_12_inst : FD1 port map( D => n5400, CP => CLK_I, Q => 
                           n_2057, QN => n3595);
   KEY_EXPAN0_reg_26_12_inst : FD1 port map( D => n5399, CP => CLK_I, Q => 
                           n_2058, QN => n3594);
   KEY_EXPAN0_reg_25_12_inst : FD1 port map( D => n5398, CP => CLK_I, Q => 
                           n_2059, QN => n3597);
   KEY_EXPAN0_reg_24_12_inst : FD1 port map( D => n5397, CP => CLK_I, Q => 
                           n_2060, QN => n3596);
   KEY_EXPAN0_reg_23_12_inst : FD1 port map( D => n5396, CP => CLK_I, Q => 
                           n_2061, QN => n3583);
   KEY_EXPAN0_reg_22_12_inst : FD1 port map( D => n5395, CP => CLK_I, Q => 
                           n_2062, QN => n3582);
   KEY_EXPAN0_reg_21_12_inst : FD1 port map( D => n5394, CP => CLK_I, Q => 
                           n_2063, QN => n3585);
   KEY_EXPAN0_reg_20_12_inst : FD1 port map( D => n5393, CP => CLK_I, Q => 
                           n_2064, QN => n3584);
   KEY_EXPAN0_reg_19_12_inst : FD1 port map( D => n5392, CP => CLK_I, Q => 
                           n_2065, QN => n3587);
   KEY_EXPAN0_reg_18_12_inst : FD1 port map( D => n5391, CP => CLK_I, Q => 
                           n_2066, QN => n3586);
   KEY_EXPAN0_reg_17_12_inst : FD1 port map( D => n5390, CP => CLK_I, Q => 
                           n_2067, QN => n3589);
   KEY_EXPAN0_reg_16_12_inst : FD1 port map( D => n5389, CP => CLK_I, Q => 
                           n_2068, QN => n3588);
   KEY_EXPAN0_reg_15_12_inst : FD1 port map( D => n5388, CP => CLK_I, Q => 
                           n_2069, QN => n3575);
   KEY_EXPAN0_reg_14_12_inst : FD1 port map( D => n5387, CP => CLK_I, Q => 
                           n_2070, QN => n3574);
   KEY_EXPAN0_reg_13_12_inst : FD1 port map( D => n5386, CP => CLK_I, Q => 
                           n_2071, QN => n3577);
   KEY_EXPAN0_reg_12_12_inst : FD1 port map( D => n5385, CP => CLK_I, Q => 
                           n_2072, QN => n3576);
   KEY_EXPAN0_reg_11_12_inst : FD1 port map( D => n5384, CP => CLK_I, Q => 
                           n_2073, QN => n3579);
   KEY_EXPAN0_reg_10_12_inst : FD1 port map( D => n5383, CP => CLK_I, Q => 
                           n_2074, QN => n3578);
   KEY_EXPAN0_reg_9_12_inst : FD1 port map( D => n5382, CP => CLK_I, Q => 
                           n_2075, QN => n3581);
   KEY_EXPAN0_reg_8_12_inst : FD1 port map( D => n5381, CP => CLK_I, Q => 
                           n_2076, QN => n3580);
   KEY_EXPAN0_reg_7_12_inst : FD1 port map( D => n5380, CP => CLK_I, Q => 
                           n_2077, QN => n3567);
   KEY_EXPAN0_reg_6_12_inst : FD1 port map( D => n5379, CP => CLK_I, Q => 
                           n_2078, QN => n3566);
   KEY_EXPAN0_reg_5_12_inst : FD1 port map( D => n5378, CP => CLK_I, Q => 
                           n_2079, QN => n3569);
   KEY_EXPAN0_reg_4_12_inst : FD1 port map( D => n5377, CP => CLK_I, Q => 
                           n_2080, QN => n3568);
   KEY_EXPAN0_reg_3_12_inst : FD1 port map( D => n5376, CP => CLK_I, Q => 
                           n_2081, QN => n3571);
   KEY_EXPAN0_reg_2_12_inst : FD1 port map( D => n5375, CP => CLK_I, Q => 
                           n_2082, QN => n3570);
   KEY_EXPAN0_reg_1_12_inst : FD1 port map( D => n5374, CP => CLK_I, Q => 
                           n_2083, QN => n3573);
   KEY_EXPAN0_reg_0_12_inst : FD1 port map( D => n5373, CP => CLK_I, Q => 
                           n_2084, QN => n3572);
   v_KEY_COL_OUT0_reg_12_inst : FD1 port map( D => n4580, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_12_port, QN => n1982);
   v_TEMP_VECTOR_reg_3_inst : FD1 port map( D => n6706, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_3_port, QN => n_2085);
   KEY_EXPAN0_reg_63_3_inst : FD1 port map( D => n4860, CP => CLK_I, Q => 
                           n_2086, QN => n3495);
   KEY_EXPAN0_reg_62_3_inst : FD1 port map( D => n4859, CP => CLK_I, Q => 
                           n_2087, QN => n3494);
   KEY_EXPAN0_reg_61_3_inst : FD1 port map( D => n4858, CP => CLK_I, Q => 
                           n_2088, QN => n3497);
   KEY_EXPAN0_reg_60_3_inst : FD1 port map( D => n4857, CP => CLK_I, Q => 
                           n_2089, QN => n3496);
   KEY_EXPAN0_reg_59_3_inst : FD1 port map( D => n4856, CP => CLK_I, Q => 
                           n_2090, QN => n3499);
   KEY_EXPAN0_reg_58_3_inst : FD1 port map( D => n4855, CP => CLK_I, Q => 
                           n_2091, QN => n3498);
   KEY_EXPAN0_reg_57_3_inst : FD1 port map( D => n4854, CP => CLK_I, Q => 
                           n_2092, QN => n3501);
   KEY_EXPAN0_reg_56_3_inst : FD1 port map( D => n4853, CP => CLK_I, Q => 
                           n_2093, QN => n3500);
   KEY_EXPAN0_reg_55_3_inst : FD1 port map( D => n4852, CP => CLK_I, Q => 
                           n_2094, QN => n3487);
   KEY_EXPAN0_reg_54_3_inst : FD1 port map( D => n4851, CP => CLK_I, Q => 
                           n_2095, QN => n3486);
   KEY_EXPAN0_reg_53_3_inst : FD1 port map( D => n4850, CP => CLK_I, Q => 
                           n_2096, QN => n3489);
   KEY_EXPAN0_reg_52_3_inst : FD1 port map( D => n4849, CP => CLK_I, Q => 
                           n_2097, QN => n3488);
   KEY_EXPAN0_reg_51_3_inst : FD1 port map( D => n4848, CP => CLK_I, Q => 
                           n_2098, QN => n3491);
   KEY_EXPAN0_reg_50_3_inst : FD1 port map( D => n4847, CP => CLK_I, Q => 
                           n_2099, QN => n3490);
   KEY_EXPAN0_reg_49_3_inst : FD1 port map( D => n4846, CP => CLK_I, Q => 
                           n_2100, QN => n3493);
   KEY_EXPAN0_reg_48_3_inst : FD1 port map( D => n4845, CP => CLK_I, Q => 
                           n_2101, QN => n3492);
   KEY_EXPAN0_reg_47_3_inst : FD1 port map( D => n4844, CP => CLK_I, Q => 
                           n_2102, QN => n3479);
   KEY_EXPAN0_reg_46_3_inst : FD1 port map( D => n4843, CP => CLK_I, Q => 
                           n_2103, QN => n3478);
   KEY_EXPAN0_reg_45_3_inst : FD1 port map( D => n4842, CP => CLK_I, Q => 
                           n_2104, QN => n3481);
   KEY_EXPAN0_reg_44_3_inst : FD1 port map( D => n4841, CP => CLK_I, Q => 
                           n_2105, QN => n3480);
   KEY_EXPAN0_reg_43_3_inst : FD1 port map( D => n4840, CP => CLK_I, Q => 
                           n_2106, QN => n3483);
   KEY_EXPAN0_reg_42_3_inst : FD1 port map( D => n4839, CP => CLK_I, Q => 
                           n_2107, QN => n3482);
   KEY_EXPAN0_reg_41_3_inst : FD1 port map( D => n4838, CP => CLK_I, Q => 
                           n_2108, QN => n3485);
   KEY_EXPAN0_reg_40_3_inst : FD1 port map( D => n4837, CP => CLK_I, Q => 
                           n_2109, QN => n3484);
   KEY_EXPAN0_reg_39_3_inst : FD1 port map( D => n4836, CP => CLK_I, Q => 
                           n_2110, QN => n3471);
   KEY_EXPAN0_reg_38_3_inst : FD1 port map( D => n4835, CP => CLK_I, Q => 
                           n_2111, QN => n3470);
   KEY_EXPAN0_reg_37_3_inst : FD1 port map( D => n4834, CP => CLK_I, Q => 
                           n_2112, QN => n3473);
   KEY_EXPAN0_reg_36_3_inst : FD1 port map( D => n4833, CP => CLK_I, Q => 
                           n_2113, QN => n3472);
   KEY_EXPAN0_reg_35_3_inst : FD1 port map( D => n4832, CP => CLK_I, Q => 
                           n_2114, QN => n3475);
   KEY_EXPAN0_reg_34_3_inst : FD1 port map( D => n4831, CP => CLK_I, Q => 
                           n_2115, QN => n3474);
   KEY_EXPAN0_reg_33_3_inst : FD1 port map( D => n4830, CP => CLK_I, Q => 
                           n_2116, QN => n3477);
   KEY_EXPAN0_reg_32_3_inst : FD1 port map( D => n4829, CP => CLK_I, Q => 
                           n_2117, QN => n3476);
   KEY_EXPAN0_reg_31_3_inst : FD1 port map( D => n4828, CP => CLK_I, Q => 
                           n_2118, QN => n3527);
   KEY_EXPAN0_reg_30_3_inst : FD1 port map( D => n4827, CP => CLK_I, Q => 
                           n_2119, QN => n3526);
   KEY_EXPAN0_reg_29_3_inst : FD1 port map( D => n4826, CP => CLK_I, Q => 
                           n_2120, QN => n3529);
   KEY_EXPAN0_reg_28_3_inst : FD1 port map( D => n4825, CP => CLK_I, Q => 
                           n_2121, QN => n3528);
   KEY_EXPAN0_reg_27_3_inst : FD1 port map( D => n4824, CP => CLK_I, Q => 
                           n_2122, QN => n3531);
   KEY_EXPAN0_reg_26_3_inst : FD1 port map( D => n4823, CP => CLK_I, Q => 
                           n_2123, QN => n3530);
   KEY_EXPAN0_reg_25_3_inst : FD1 port map( D => n4822, CP => CLK_I, Q => 
                           n_2124, QN => n3533);
   KEY_EXPAN0_reg_24_3_inst : FD1 port map( D => n4821, CP => CLK_I, Q => 
                           n_2125, QN => n3532);
   KEY_EXPAN0_reg_23_3_inst : FD1 port map( D => n4820, CP => CLK_I, Q => 
                           n_2126, QN => n3519);
   KEY_EXPAN0_reg_22_3_inst : FD1 port map( D => n4819, CP => CLK_I, Q => 
                           n_2127, QN => n3518);
   KEY_EXPAN0_reg_21_3_inst : FD1 port map( D => n4818, CP => CLK_I, Q => 
                           n_2128, QN => n3521);
   KEY_EXPAN0_reg_20_3_inst : FD1 port map( D => n4817, CP => CLK_I, Q => 
                           n_2129, QN => n3520);
   KEY_EXPAN0_reg_19_3_inst : FD1 port map( D => n4816, CP => CLK_I, Q => 
                           n_2130, QN => n3523);
   KEY_EXPAN0_reg_18_3_inst : FD1 port map( D => n4815, CP => CLK_I, Q => 
                           n_2131, QN => n3522);
   KEY_EXPAN0_reg_17_3_inst : FD1 port map( D => n4814, CP => CLK_I, Q => 
                           n_2132, QN => n3525);
   KEY_EXPAN0_reg_16_3_inst : FD1 port map( D => n4813, CP => CLK_I, Q => 
                           n_2133, QN => n3524);
   KEY_EXPAN0_reg_15_3_inst : FD1 port map( D => n4812, CP => CLK_I, Q => 
                           n_2134, QN => n3511);
   KEY_EXPAN0_reg_14_3_inst : FD1 port map( D => n4811, CP => CLK_I, Q => 
                           n_2135, QN => n3510);
   KEY_EXPAN0_reg_13_3_inst : FD1 port map( D => n4810, CP => CLK_I, Q => 
                           n_2136, QN => n3513);
   KEY_EXPAN0_reg_12_3_inst : FD1 port map( D => n4809, CP => CLK_I, Q => 
                           n_2137, QN => n3512);
   KEY_EXPAN0_reg_11_3_inst : FD1 port map( D => n4808, CP => CLK_I, Q => 
                           n_2138, QN => n3515);
   KEY_EXPAN0_reg_10_3_inst : FD1 port map( D => n4807, CP => CLK_I, Q => 
                           n_2139, QN => n3514);
   KEY_EXPAN0_reg_9_3_inst : FD1 port map( D => n4806, CP => CLK_I, Q => n_2140
                           , QN => n3517);
   KEY_EXPAN0_reg_8_3_inst : FD1 port map( D => n4805, CP => CLK_I, Q => n_2141
                           , QN => n3516);
   KEY_EXPAN0_reg_7_3_inst : FD1 port map( D => n4804, CP => CLK_I, Q => n_2142
                           , QN => n3503);
   KEY_EXPAN0_reg_6_3_inst : FD1 port map( D => n4803, CP => CLK_I, Q => n_2143
                           , QN => n3502);
   KEY_EXPAN0_reg_5_3_inst : FD1 port map( D => n4802, CP => CLK_I, Q => n_2144
                           , QN => n3505);
   KEY_EXPAN0_reg_4_3_inst : FD1 port map( D => n4801, CP => CLK_I, Q => n_2145
                           , QN => n3504);
   KEY_EXPAN0_reg_3_3_inst : FD1 port map( D => n4800, CP => CLK_I, Q => n_2146
                           , QN => n3507);
   KEY_EXPAN0_reg_2_3_inst : FD1 port map( D => n4799, CP => CLK_I, Q => n_2147
                           , QN => n3506);
   KEY_EXPAN0_reg_1_3_inst : FD1 port map( D => n4798, CP => CLK_I, Q => n_2148
                           , QN => n3509);
   KEY_EXPAN0_reg_0_3_inst : FD1 port map( D => n4797, CP => CLK_I, Q => n_2149
                           , QN => n3508);
   v_KEY_COL_OUT0_reg_3_inst : FD1 port map( D => n4579, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_3_port, QN => n2001);
   v_TEMP_VECTOR_reg_27_inst : FD1 port map( D => n6682, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_27_port, QN => n_2150);
   KEY_EXPAN0_reg_63_27_inst : FD1 port map( D => n6396, CP => CLK_I, Q => 
                           n_2151, QN => n3431);
   KEY_EXPAN0_reg_62_27_inst : FD1 port map( D => n6395, CP => CLK_I, Q => 
                           n_2152, QN => n3430);
   KEY_EXPAN0_reg_61_27_inst : FD1 port map( D => n6394, CP => CLK_I, Q => 
                           n_2153, QN => n3433);
   KEY_EXPAN0_reg_60_27_inst : FD1 port map( D => n6393, CP => CLK_I, Q => 
                           n_2154, QN => n3432);
   KEY_EXPAN0_reg_59_27_inst : FD1 port map( D => n6392, CP => CLK_I, Q => 
                           n_2155, QN => n3435);
   KEY_EXPAN0_reg_58_27_inst : FD1 port map( D => n6391, CP => CLK_I, Q => 
                           n_2156, QN => n3434);
   KEY_EXPAN0_reg_57_27_inst : FD1 port map( D => n6390, CP => CLK_I, Q => 
                           n_2157, QN => n3437);
   KEY_EXPAN0_reg_56_27_inst : FD1 port map( D => n6389, CP => CLK_I, Q => 
                           n_2158, QN => n3436);
   KEY_EXPAN0_reg_55_27_inst : FD1 port map( D => n6388, CP => CLK_I, Q => 
                           n_2159, QN => n3423);
   KEY_EXPAN0_reg_54_27_inst : FD1 port map( D => n6387, CP => CLK_I, Q => 
                           n_2160, QN => n3422);
   KEY_EXPAN0_reg_53_27_inst : FD1 port map( D => n6386, CP => CLK_I, Q => 
                           n_2161, QN => n3425);
   KEY_EXPAN0_reg_52_27_inst : FD1 port map( D => n6385, CP => CLK_I, Q => 
                           n_2162, QN => n3424);
   KEY_EXPAN0_reg_51_27_inst : FD1 port map( D => n6384, CP => CLK_I, Q => 
                           n_2163, QN => n3427);
   KEY_EXPAN0_reg_50_27_inst : FD1 port map( D => n6383, CP => CLK_I, Q => 
                           n_2164, QN => n3426);
   KEY_EXPAN0_reg_49_27_inst : FD1 port map( D => n6382, CP => CLK_I, Q => 
                           n_2165, QN => n3429);
   KEY_EXPAN0_reg_48_27_inst : FD1 port map( D => n6381, CP => CLK_I, Q => 
                           n_2166, QN => n3428);
   KEY_EXPAN0_reg_47_27_inst : FD1 port map( D => n6380, CP => CLK_I, Q => 
                           n_2167, QN => n3415);
   KEY_EXPAN0_reg_46_27_inst : FD1 port map( D => n6379, CP => CLK_I, Q => 
                           n_2168, QN => n3414);
   KEY_EXPAN0_reg_45_27_inst : FD1 port map( D => n6378, CP => CLK_I, Q => 
                           n_2169, QN => n3417);
   KEY_EXPAN0_reg_44_27_inst : FD1 port map( D => n6377, CP => CLK_I, Q => 
                           n_2170, QN => n3416);
   KEY_EXPAN0_reg_43_27_inst : FD1 port map( D => n6376, CP => CLK_I, Q => 
                           n_2171, QN => n3419);
   KEY_EXPAN0_reg_42_27_inst : FD1 port map( D => n6375, CP => CLK_I, Q => 
                           n_2172, QN => n3418);
   KEY_EXPAN0_reg_41_27_inst : FD1 port map( D => n6374, CP => CLK_I, Q => 
                           n_2173, QN => n3421);
   KEY_EXPAN0_reg_40_27_inst : FD1 port map( D => n6373, CP => CLK_I, Q => 
                           n_2174, QN => n3420);
   KEY_EXPAN0_reg_39_27_inst : FD1 port map( D => n6372, CP => CLK_I, Q => 
                           n_2175, QN => n3407);
   KEY_EXPAN0_reg_38_27_inst : FD1 port map( D => n6371, CP => CLK_I, Q => 
                           n_2176, QN => n3406);
   KEY_EXPAN0_reg_37_27_inst : FD1 port map( D => n6370, CP => CLK_I, Q => 
                           n_2177, QN => n3409);
   KEY_EXPAN0_reg_36_27_inst : FD1 port map( D => n6369, CP => CLK_I, Q => 
                           n_2178, QN => n3408);
   KEY_EXPAN0_reg_35_27_inst : FD1 port map( D => n6368, CP => CLK_I, Q => 
                           n_2179, QN => n3411);
   KEY_EXPAN0_reg_34_27_inst : FD1 port map( D => n6367, CP => CLK_I, Q => 
                           n_2180, QN => n3410);
   KEY_EXPAN0_reg_33_27_inst : FD1 port map( D => n6366, CP => CLK_I, Q => 
                           n_2181, QN => n3413);
   KEY_EXPAN0_reg_32_27_inst : FD1 port map( D => n6365, CP => CLK_I, Q => 
                           n_2182, QN => n3412);
   KEY_EXPAN0_reg_31_27_inst : FD1 port map( D => n6364, CP => CLK_I, Q => 
                           n_2183, QN => n3463);
   KEY_EXPAN0_reg_30_27_inst : FD1 port map( D => n6363, CP => CLK_I, Q => 
                           n_2184, QN => n3462);
   KEY_EXPAN0_reg_29_27_inst : FD1 port map( D => n6362, CP => CLK_I, Q => 
                           n_2185, QN => n3465);
   KEY_EXPAN0_reg_28_27_inst : FD1 port map( D => n6361, CP => CLK_I, Q => 
                           n_2186, QN => n3464);
   KEY_EXPAN0_reg_27_27_inst : FD1 port map( D => n6360, CP => CLK_I, Q => 
                           n_2187, QN => n3467);
   KEY_EXPAN0_reg_26_27_inst : FD1 port map( D => n6359, CP => CLK_I, Q => 
                           n_2188, QN => n3466);
   KEY_EXPAN0_reg_25_27_inst : FD1 port map( D => n6358, CP => CLK_I, Q => 
                           n_2189, QN => n3469);
   KEY_EXPAN0_reg_24_27_inst : FD1 port map( D => n6357, CP => CLK_I, Q => 
                           n_2190, QN => n3468);
   KEY_EXPAN0_reg_23_27_inst : FD1 port map( D => n6356, CP => CLK_I, Q => 
                           n_2191, QN => n3455);
   KEY_EXPAN0_reg_22_27_inst : FD1 port map( D => n6355, CP => CLK_I, Q => 
                           n_2192, QN => n3454);
   KEY_EXPAN0_reg_21_27_inst : FD1 port map( D => n6354, CP => CLK_I, Q => 
                           n_2193, QN => n3457);
   KEY_EXPAN0_reg_20_27_inst : FD1 port map( D => n6353, CP => CLK_I, Q => 
                           n_2194, QN => n3456);
   KEY_EXPAN0_reg_19_27_inst : FD1 port map( D => n6352, CP => CLK_I, Q => 
                           n_2195, QN => n3459);
   KEY_EXPAN0_reg_18_27_inst : FD1 port map( D => n6351, CP => CLK_I, Q => 
                           n_2196, QN => n3458);
   KEY_EXPAN0_reg_17_27_inst : FD1 port map( D => n6350, CP => CLK_I, Q => 
                           n_2197, QN => n3461);
   KEY_EXPAN0_reg_16_27_inst : FD1 port map( D => n6349, CP => CLK_I, Q => 
                           n_2198, QN => n3460);
   KEY_EXPAN0_reg_15_27_inst : FD1 port map( D => n6348, CP => CLK_I, Q => 
                           n_2199, QN => n3447);
   KEY_EXPAN0_reg_14_27_inst : FD1 port map( D => n6347, CP => CLK_I, Q => 
                           n_2200, QN => n3446);
   KEY_EXPAN0_reg_13_27_inst : FD1 port map( D => n6346, CP => CLK_I, Q => 
                           n_2201, QN => n3449);
   KEY_EXPAN0_reg_12_27_inst : FD1 port map( D => n6345, CP => CLK_I, Q => 
                           n_2202, QN => n3448);
   KEY_EXPAN0_reg_11_27_inst : FD1 port map( D => n6344, CP => CLK_I, Q => 
                           n_2203, QN => n3451);
   KEY_EXPAN0_reg_10_27_inst : FD1 port map( D => n6343, CP => CLK_I, Q => 
                           n_2204, QN => n3450);
   KEY_EXPAN0_reg_9_27_inst : FD1 port map( D => n6342, CP => CLK_I, Q => 
                           n_2205, QN => n3453);
   KEY_EXPAN0_reg_8_27_inst : FD1 port map( D => n6341, CP => CLK_I, Q => 
                           n_2206, QN => n3452);
   KEY_EXPAN0_reg_7_27_inst : FD1 port map( D => n6340, CP => CLK_I, Q => 
                           n_2207, QN => n3439);
   KEY_EXPAN0_reg_6_27_inst : FD1 port map( D => n6339, CP => CLK_I, Q => 
                           n_2208, QN => n3438);
   KEY_EXPAN0_reg_5_27_inst : FD1 port map( D => n6338, CP => CLK_I, Q => 
                           n_2209, QN => n3441);
   KEY_EXPAN0_reg_4_27_inst : FD1 port map( D => n6337, CP => CLK_I, Q => 
                           n_2210, QN => n3440);
   KEY_EXPAN0_reg_3_27_inst : FD1 port map( D => n6336, CP => CLK_I, Q => 
                           n_2211, QN => n3443);
   KEY_EXPAN0_reg_2_27_inst : FD1 port map( D => n6335, CP => CLK_I, Q => 
                           n_2212, QN => n3442);
   KEY_EXPAN0_reg_1_27_inst : FD1 port map( D => n6334, CP => CLK_I, Q => 
                           n_2213, QN => n3445);
   KEY_EXPAN0_reg_0_27_inst : FD1 port map( D => n6333, CP => CLK_I, Q => 
                           n_2214, QN => n3444);
   v_KEY_COL_OUT0_reg_27_inst : FD1 port map( D => n4578, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_27_port, QN => n1868);
   v_TEMP_VECTOR_reg_19_inst : FD1 port map( D => n6690, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_19_port, QN => n_2215);
   KEY_EXPAN0_reg_63_19_inst : FD1 port map( D => n5884, CP => CLK_I, Q => 
                           n_2216, QN => n3367);
   KEY_EXPAN0_reg_62_19_inst : FD1 port map( D => n5883, CP => CLK_I, Q => 
                           n_2217, QN => n3366);
   KEY_EXPAN0_reg_61_19_inst : FD1 port map( D => n5882, CP => CLK_I, Q => 
                           n_2218, QN => n3369);
   KEY_EXPAN0_reg_60_19_inst : FD1 port map( D => n5881, CP => CLK_I, Q => 
                           n_2219, QN => n3368);
   KEY_EXPAN0_reg_59_19_inst : FD1 port map( D => n5880, CP => CLK_I, Q => 
                           n_2220, QN => n3371);
   KEY_EXPAN0_reg_58_19_inst : FD1 port map( D => n5879, CP => CLK_I, Q => 
                           n_2221, QN => n3370);
   KEY_EXPAN0_reg_57_19_inst : FD1 port map( D => n5878, CP => CLK_I, Q => 
                           n_2222, QN => n3373);
   KEY_EXPAN0_reg_56_19_inst : FD1 port map( D => n5877, CP => CLK_I, Q => 
                           n_2223, QN => n3372);
   KEY_EXPAN0_reg_55_19_inst : FD1 port map( D => n5876, CP => CLK_I, Q => 
                           n_2224, QN => n3359);
   KEY_EXPAN0_reg_54_19_inst : FD1 port map( D => n5875, CP => CLK_I, Q => 
                           n_2225, QN => n3358);
   KEY_EXPAN0_reg_53_19_inst : FD1 port map( D => n5874, CP => CLK_I, Q => 
                           n_2226, QN => n3361);
   KEY_EXPAN0_reg_52_19_inst : FD1 port map( D => n5873, CP => CLK_I, Q => 
                           n_2227, QN => n3360);
   KEY_EXPAN0_reg_51_19_inst : FD1 port map( D => n5872, CP => CLK_I, Q => 
                           n_2228, QN => n3363);
   KEY_EXPAN0_reg_50_19_inst : FD1 port map( D => n5871, CP => CLK_I, Q => 
                           n_2229, QN => n3362);
   KEY_EXPAN0_reg_49_19_inst : FD1 port map( D => n5870, CP => CLK_I, Q => 
                           n_2230, QN => n3365);
   KEY_EXPAN0_reg_48_19_inst : FD1 port map( D => n5869, CP => CLK_I, Q => 
                           n_2231, QN => n3364);
   KEY_EXPAN0_reg_47_19_inst : FD1 port map( D => n5868, CP => CLK_I, Q => 
                           n_2232, QN => n3351);
   KEY_EXPAN0_reg_46_19_inst : FD1 port map( D => n5867, CP => CLK_I, Q => 
                           n_2233, QN => n3350);
   KEY_EXPAN0_reg_45_19_inst : FD1 port map( D => n5866, CP => CLK_I, Q => 
                           n_2234, QN => n3353);
   KEY_EXPAN0_reg_44_19_inst : FD1 port map( D => n5865, CP => CLK_I, Q => 
                           n_2235, QN => n3352);
   KEY_EXPAN0_reg_43_19_inst : FD1 port map( D => n5864, CP => CLK_I, Q => 
                           n_2236, QN => n3355);
   KEY_EXPAN0_reg_42_19_inst : FD1 port map( D => n5863, CP => CLK_I, Q => 
                           n_2237, QN => n3354);
   KEY_EXPAN0_reg_41_19_inst : FD1 port map( D => n5862, CP => CLK_I, Q => 
                           n_2238, QN => n3357);
   KEY_EXPAN0_reg_40_19_inst : FD1 port map( D => n5861, CP => CLK_I, Q => 
                           n_2239, QN => n3356);
   KEY_EXPAN0_reg_39_19_inst : FD1 port map( D => n5860, CP => CLK_I, Q => 
                           n_2240, QN => n3343);
   KEY_EXPAN0_reg_38_19_inst : FD1 port map( D => n5859, CP => CLK_I, Q => 
                           n_2241, QN => n3342);
   KEY_EXPAN0_reg_37_19_inst : FD1 port map( D => n5858, CP => CLK_I, Q => 
                           n_2242, QN => n3345);
   KEY_EXPAN0_reg_36_19_inst : FD1 port map( D => n5857, CP => CLK_I, Q => 
                           n_2243, QN => n3344);
   KEY_EXPAN0_reg_35_19_inst : FD1 port map( D => n5856, CP => CLK_I, Q => 
                           n_2244, QN => n3347);
   KEY_EXPAN0_reg_34_19_inst : FD1 port map( D => n5855, CP => CLK_I, Q => 
                           n_2245, QN => n3346);
   KEY_EXPAN0_reg_33_19_inst : FD1 port map( D => n5854, CP => CLK_I, Q => 
                           n_2246, QN => n3349);
   KEY_EXPAN0_reg_32_19_inst : FD1 port map( D => n5853, CP => CLK_I, Q => 
                           n_2247, QN => n3348);
   KEY_EXPAN0_reg_31_19_inst : FD1 port map( D => n5852, CP => CLK_I, Q => 
                           n_2248, QN => n3399);
   KEY_EXPAN0_reg_30_19_inst : FD1 port map( D => n5851, CP => CLK_I, Q => 
                           n_2249, QN => n3398);
   KEY_EXPAN0_reg_29_19_inst : FD1 port map( D => n5850, CP => CLK_I, Q => 
                           n_2250, QN => n3401);
   KEY_EXPAN0_reg_28_19_inst : FD1 port map( D => n5849, CP => CLK_I, Q => 
                           n_2251, QN => n3400);
   KEY_EXPAN0_reg_27_19_inst : FD1 port map( D => n5848, CP => CLK_I, Q => 
                           n_2252, QN => n3403);
   KEY_EXPAN0_reg_26_19_inst : FD1 port map( D => n5847, CP => CLK_I, Q => 
                           n_2253, QN => n3402);
   KEY_EXPAN0_reg_25_19_inst : FD1 port map( D => n5846, CP => CLK_I, Q => 
                           n_2254, QN => n3405);
   KEY_EXPAN0_reg_24_19_inst : FD1 port map( D => n5845, CP => CLK_I, Q => 
                           n_2255, QN => n3404);
   KEY_EXPAN0_reg_23_19_inst : FD1 port map( D => n5844, CP => CLK_I, Q => 
                           n_2256, QN => n3391);
   KEY_EXPAN0_reg_22_19_inst : FD1 port map( D => n5843, CP => CLK_I, Q => 
                           n_2257, QN => n3390);
   KEY_EXPAN0_reg_21_19_inst : FD1 port map( D => n5842, CP => CLK_I, Q => 
                           n_2258, QN => n3393);
   KEY_EXPAN0_reg_20_19_inst : FD1 port map( D => n5841, CP => CLK_I, Q => 
                           n_2259, QN => n3392);
   KEY_EXPAN0_reg_19_19_inst : FD1 port map( D => n5840, CP => CLK_I, Q => 
                           n_2260, QN => n3395);
   KEY_EXPAN0_reg_18_19_inst : FD1 port map( D => n5839, CP => CLK_I, Q => 
                           n_2261, QN => n3394);
   KEY_EXPAN0_reg_17_19_inst : FD1 port map( D => n5838, CP => CLK_I, Q => 
                           n_2262, QN => n3397);
   KEY_EXPAN0_reg_16_19_inst : FD1 port map( D => n5837, CP => CLK_I, Q => 
                           n_2263, QN => n3396);
   KEY_EXPAN0_reg_15_19_inst : FD1 port map( D => n5836, CP => CLK_I, Q => 
                           n_2264, QN => n3383);
   KEY_EXPAN0_reg_14_19_inst : FD1 port map( D => n5835, CP => CLK_I, Q => 
                           n_2265, QN => n3382);
   KEY_EXPAN0_reg_13_19_inst : FD1 port map( D => n5834, CP => CLK_I, Q => 
                           n_2266, QN => n3385);
   KEY_EXPAN0_reg_12_19_inst : FD1 port map( D => n5833, CP => CLK_I, Q => 
                           n_2267, QN => n3384);
   KEY_EXPAN0_reg_11_19_inst : FD1 port map( D => n5832, CP => CLK_I, Q => 
                           n_2268, QN => n3387);
   KEY_EXPAN0_reg_10_19_inst : FD1 port map( D => n5831, CP => CLK_I, Q => 
                           n_2269, QN => n3386);
   KEY_EXPAN0_reg_9_19_inst : FD1 port map( D => n5830, CP => CLK_I, Q => 
                           n_2270, QN => n3389);
   KEY_EXPAN0_reg_8_19_inst : FD1 port map( D => n5829, CP => CLK_I, Q => 
                           n_2271, QN => n3388);
   KEY_EXPAN0_reg_7_19_inst : FD1 port map( D => n5828, CP => CLK_I, Q => 
                           n_2272, QN => n3375);
   KEY_EXPAN0_reg_6_19_inst : FD1 port map( D => n5827, CP => CLK_I, Q => 
                           n_2273, QN => n3374);
   KEY_EXPAN0_reg_5_19_inst : FD1 port map( D => n5826, CP => CLK_I, Q => 
                           n_2274, QN => n3377);
   KEY_EXPAN0_reg_4_19_inst : FD1 port map( D => n5825, CP => CLK_I, Q => 
                           n_2275, QN => n3376);
   KEY_EXPAN0_reg_3_19_inst : FD1 port map( D => n5824, CP => CLK_I, Q => 
                           n_2276, QN => n3379);
   KEY_EXPAN0_reg_2_19_inst : FD1 port map( D => n5823, CP => CLK_I, Q => 
                           n_2277, QN => n3378);
   KEY_EXPAN0_reg_1_19_inst : FD1 port map( D => n5822, CP => CLK_I, Q => 
                           n_2278, QN => n3381);
   KEY_EXPAN0_reg_0_19_inst : FD1 port map( D => n5821, CP => CLK_I, Q => 
                           n_2279, QN => n3380);
   v_KEY_COL_OUT0_reg_19_inst : FD1 port map( D => n4577, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_19_port, QN => n1962);
   v_TEMP_VECTOR_reg_11_inst : FD1 port map( D => n6698, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_11_port, QN => n_2280);
   KEY_EXPAN0_reg_63_11_inst : FD1 port map( D => n5372, CP => CLK_I, Q => 
                           n_2281, QN => n3303);
   KEY_EXPAN0_reg_62_11_inst : FD1 port map( D => n5371, CP => CLK_I, Q => 
                           n_2282, QN => n3302);
   KEY_EXPAN0_reg_61_11_inst : FD1 port map( D => n5370, CP => CLK_I, Q => 
                           n_2283, QN => n3305);
   KEY_EXPAN0_reg_60_11_inst : FD1 port map( D => n5369, CP => CLK_I, Q => 
                           n_2284, QN => n3304);
   KEY_EXPAN0_reg_59_11_inst : FD1 port map( D => n5368, CP => CLK_I, Q => 
                           n_2285, QN => n3307);
   KEY_EXPAN0_reg_58_11_inst : FD1 port map( D => n5367, CP => CLK_I, Q => 
                           n_2286, QN => n3306);
   KEY_EXPAN0_reg_57_11_inst : FD1 port map( D => n5366, CP => CLK_I, Q => 
                           n_2287, QN => n3309);
   KEY_EXPAN0_reg_56_11_inst : FD1 port map( D => n5365, CP => CLK_I, Q => 
                           n_2288, QN => n3308);
   KEY_EXPAN0_reg_55_11_inst : FD1 port map( D => n5364, CP => CLK_I, Q => 
                           n_2289, QN => n3295);
   KEY_EXPAN0_reg_54_11_inst : FD1 port map( D => n5363, CP => CLK_I, Q => 
                           n_2290, QN => n3294);
   KEY_EXPAN0_reg_53_11_inst : FD1 port map( D => n5362, CP => CLK_I, Q => 
                           n_2291, QN => n3297);
   KEY_EXPAN0_reg_52_11_inst : FD1 port map( D => n5361, CP => CLK_I, Q => 
                           n_2292, QN => n3296);
   KEY_EXPAN0_reg_51_11_inst : FD1 port map( D => n5360, CP => CLK_I, Q => 
                           n_2293, QN => n3299);
   KEY_EXPAN0_reg_50_11_inst : FD1 port map( D => n5359, CP => CLK_I, Q => 
                           n_2294, QN => n3298);
   KEY_EXPAN0_reg_49_11_inst : FD1 port map( D => n5358, CP => CLK_I, Q => 
                           n_2295, QN => n3301);
   KEY_EXPAN0_reg_48_11_inst : FD1 port map( D => n5357, CP => CLK_I, Q => 
                           n_2296, QN => n3300);
   KEY_EXPAN0_reg_47_11_inst : FD1 port map( D => n5356, CP => CLK_I, Q => 
                           n_2297, QN => n3287);
   KEY_EXPAN0_reg_46_11_inst : FD1 port map( D => n5355, CP => CLK_I, Q => 
                           n_2298, QN => n3286);
   KEY_EXPAN0_reg_45_11_inst : FD1 port map( D => n5354, CP => CLK_I, Q => 
                           n_2299, QN => n3289);
   KEY_EXPAN0_reg_44_11_inst : FD1 port map( D => n5353, CP => CLK_I, Q => 
                           n_2300, QN => n3288);
   KEY_EXPAN0_reg_43_11_inst : FD1 port map( D => n5352, CP => CLK_I, Q => 
                           n_2301, QN => n3291);
   KEY_EXPAN0_reg_42_11_inst : FD1 port map( D => n5351, CP => CLK_I, Q => 
                           n_2302, QN => n3290);
   KEY_EXPAN0_reg_41_11_inst : FD1 port map( D => n5350, CP => CLK_I, Q => 
                           n_2303, QN => n3293);
   KEY_EXPAN0_reg_40_11_inst : FD1 port map( D => n5349, CP => CLK_I, Q => 
                           n_2304, QN => n3292);
   KEY_EXPAN0_reg_39_11_inst : FD1 port map( D => n5348, CP => CLK_I, Q => 
                           n_2305, QN => n3279);
   KEY_EXPAN0_reg_38_11_inst : FD1 port map( D => n5347, CP => CLK_I, Q => 
                           n_2306, QN => n3278);
   KEY_EXPAN0_reg_37_11_inst : FD1 port map( D => n5346, CP => CLK_I, Q => 
                           n_2307, QN => n3281);
   KEY_EXPAN0_reg_36_11_inst : FD1 port map( D => n5345, CP => CLK_I, Q => 
                           n_2308, QN => n3280);
   KEY_EXPAN0_reg_35_11_inst : FD1 port map( D => n5344, CP => CLK_I, Q => 
                           n_2309, QN => n3283);
   KEY_EXPAN0_reg_34_11_inst : FD1 port map( D => n5343, CP => CLK_I, Q => 
                           n_2310, QN => n3282);
   KEY_EXPAN0_reg_33_11_inst : FD1 port map( D => n5342, CP => CLK_I, Q => 
                           n_2311, QN => n3285);
   KEY_EXPAN0_reg_32_11_inst : FD1 port map( D => n5341, CP => CLK_I, Q => 
                           n_2312, QN => n3284);
   KEY_EXPAN0_reg_31_11_inst : FD1 port map( D => n5340, CP => CLK_I, Q => 
                           n_2313, QN => n3335);
   KEY_EXPAN0_reg_30_11_inst : FD1 port map( D => n5339, CP => CLK_I, Q => 
                           n_2314, QN => n3334);
   KEY_EXPAN0_reg_29_11_inst : FD1 port map( D => n5338, CP => CLK_I, Q => 
                           n_2315, QN => n3337);
   KEY_EXPAN0_reg_28_11_inst : FD1 port map( D => n5337, CP => CLK_I, Q => 
                           n_2316, QN => n3336);
   KEY_EXPAN0_reg_27_11_inst : FD1 port map( D => n5336, CP => CLK_I, Q => 
                           n_2317, QN => n3339);
   KEY_EXPAN0_reg_26_11_inst : FD1 port map( D => n5335, CP => CLK_I, Q => 
                           n_2318, QN => n3338);
   KEY_EXPAN0_reg_25_11_inst : FD1 port map( D => n5334, CP => CLK_I, Q => 
                           n_2319, QN => n3341);
   KEY_EXPAN0_reg_24_11_inst : FD1 port map( D => n5333, CP => CLK_I, Q => 
                           n_2320, QN => n3340);
   KEY_EXPAN0_reg_23_11_inst : FD1 port map( D => n5332, CP => CLK_I, Q => 
                           n_2321, QN => n3327);
   KEY_EXPAN0_reg_22_11_inst : FD1 port map( D => n5331, CP => CLK_I, Q => 
                           n_2322, QN => n3326);
   KEY_EXPAN0_reg_21_11_inst : FD1 port map( D => n5330, CP => CLK_I, Q => 
                           n_2323, QN => n3329);
   KEY_EXPAN0_reg_20_11_inst : FD1 port map( D => n5329, CP => CLK_I, Q => 
                           n_2324, QN => n3328);
   KEY_EXPAN0_reg_19_11_inst : FD1 port map( D => n5328, CP => CLK_I, Q => 
                           n_2325, QN => n3331);
   KEY_EXPAN0_reg_18_11_inst : FD1 port map( D => n5327, CP => CLK_I, Q => 
                           n_2326, QN => n3330);
   KEY_EXPAN0_reg_17_11_inst : FD1 port map( D => n5326, CP => CLK_I, Q => 
                           n_2327, QN => n3333);
   KEY_EXPAN0_reg_16_11_inst : FD1 port map( D => n5325, CP => CLK_I, Q => 
                           n_2328, QN => n3332);
   KEY_EXPAN0_reg_15_11_inst : FD1 port map( D => n5324, CP => CLK_I, Q => 
                           n_2329, QN => n3319);
   KEY_EXPAN0_reg_14_11_inst : FD1 port map( D => n5323, CP => CLK_I, Q => 
                           n_2330, QN => n3318);
   KEY_EXPAN0_reg_13_11_inst : FD1 port map( D => n5322, CP => CLK_I, Q => 
                           n_2331, QN => n3321);
   KEY_EXPAN0_reg_12_11_inst : FD1 port map( D => n5321, CP => CLK_I, Q => 
                           n_2332, QN => n3320);
   KEY_EXPAN0_reg_11_11_inst : FD1 port map( D => n5320, CP => CLK_I, Q => 
                           n_2333, QN => n3323);
   KEY_EXPAN0_reg_10_11_inst : FD1 port map( D => n5319, CP => CLK_I, Q => 
                           n_2334, QN => n3322);
   KEY_EXPAN0_reg_9_11_inst : FD1 port map( D => n5318, CP => CLK_I, Q => 
                           n_2335, QN => n3325);
   KEY_EXPAN0_reg_8_11_inst : FD1 port map( D => n5317, CP => CLK_I, Q => 
                           n_2336, QN => n3324);
   KEY_EXPAN0_reg_7_11_inst : FD1 port map( D => n5316, CP => CLK_I, Q => 
                           n_2337, QN => n3311);
   KEY_EXPAN0_reg_6_11_inst : FD1 port map( D => n5315, CP => CLK_I, Q => 
                           n_2338, QN => n3310);
   KEY_EXPAN0_reg_5_11_inst : FD1 port map( D => n5314, CP => CLK_I, Q => 
                           n_2339, QN => n3313);
   KEY_EXPAN0_reg_4_11_inst : FD1 port map( D => n5313, CP => CLK_I, Q => 
                           n_2340, QN => n3312);
   KEY_EXPAN0_reg_3_11_inst : FD1 port map( D => n5312, CP => CLK_I, Q => 
                           n_2341, QN => n3315);
   KEY_EXPAN0_reg_2_11_inst : FD1 port map( D => n5311, CP => CLK_I, Q => 
                           n_2342, QN => n3314);
   KEY_EXPAN0_reg_1_11_inst : FD1 port map( D => n5310, CP => CLK_I, Q => 
                           n_2343, QN => n3317);
   KEY_EXPAN0_reg_0_11_inst : FD1 port map( D => n5309, CP => CLK_I, Q => 
                           n_2344, QN => n3316);
   v_KEY_COL_OUT0_reg_11_inst : FD1 port map( D => n4576, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_11_port, QN => n1872);
   v_TEMP_VECTOR_reg_2_inst : FD1 port map( D => n6707, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_2_port, QN => n_2345);
   KEY_EXPAN0_reg_63_2_inst : FD1 port map( D => n4796, CP => CLK_I, Q => 
                           n_2346, QN => n3239);
   KEY_EXPAN0_reg_62_2_inst : FD1 port map( D => n4795, CP => CLK_I, Q => 
                           n_2347, QN => n3238);
   KEY_EXPAN0_reg_61_2_inst : FD1 port map( D => n4794, CP => CLK_I, Q => 
                           n_2348, QN => n3241);
   KEY_EXPAN0_reg_60_2_inst : FD1 port map( D => n4793, CP => CLK_I, Q => 
                           n_2349, QN => n3240);
   KEY_EXPAN0_reg_59_2_inst : FD1 port map( D => n4792, CP => CLK_I, Q => 
                           n_2350, QN => n3243);
   KEY_EXPAN0_reg_58_2_inst : FD1 port map( D => n4791, CP => CLK_I, Q => 
                           n_2351, QN => n3242);
   KEY_EXPAN0_reg_57_2_inst : FD1 port map( D => n4790, CP => CLK_I, Q => 
                           n_2352, QN => n3245);
   KEY_EXPAN0_reg_56_2_inst : FD1 port map( D => n4789, CP => CLK_I, Q => 
                           n_2353, QN => n3244);
   KEY_EXPAN0_reg_55_2_inst : FD1 port map( D => n4788, CP => CLK_I, Q => 
                           n_2354, QN => n3231);
   KEY_EXPAN0_reg_54_2_inst : FD1 port map( D => n4787, CP => CLK_I, Q => 
                           n_2355, QN => n3230);
   KEY_EXPAN0_reg_53_2_inst : FD1 port map( D => n4786, CP => CLK_I, Q => 
                           n_2356, QN => n3233);
   KEY_EXPAN0_reg_52_2_inst : FD1 port map( D => n4785, CP => CLK_I, Q => 
                           n_2357, QN => n3232);
   KEY_EXPAN0_reg_51_2_inst : FD1 port map( D => n4784, CP => CLK_I, Q => 
                           n_2358, QN => n3235);
   KEY_EXPAN0_reg_50_2_inst : FD1 port map( D => n4783, CP => CLK_I, Q => 
                           n_2359, QN => n3234);
   KEY_EXPAN0_reg_49_2_inst : FD1 port map( D => n4782, CP => CLK_I, Q => 
                           n_2360, QN => n3237);
   KEY_EXPAN0_reg_48_2_inst : FD1 port map( D => n4781, CP => CLK_I, Q => 
                           n_2361, QN => n3236);
   KEY_EXPAN0_reg_47_2_inst : FD1 port map( D => n4780, CP => CLK_I, Q => 
                           n_2362, QN => n3223);
   KEY_EXPAN0_reg_46_2_inst : FD1 port map( D => n4779, CP => CLK_I, Q => 
                           n_2363, QN => n3222);
   KEY_EXPAN0_reg_45_2_inst : FD1 port map( D => n4778, CP => CLK_I, Q => 
                           n_2364, QN => n3225);
   KEY_EXPAN0_reg_44_2_inst : FD1 port map( D => n4777, CP => CLK_I, Q => 
                           n_2365, QN => n3224);
   KEY_EXPAN0_reg_43_2_inst : FD1 port map( D => n4776, CP => CLK_I, Q => 
                           n_2366, QN => n3227);
   KEY_EXPAN0_reg_42_2_inst : FD1 port map( D => n4775, CP => CLK_I, Q => 
                           n_2367, QN => n3226);
   KEY_EXPAN0_reg_41_2_inst : FD1 port map( D => n4774, CP => CLK_I, Q => 
                           n_2368, QN => n3229);
   KEY_EXPAN0_reg_40_2_inst : FD1 port map( D => n4773, CP => CLK_I, Q => 
                           n_2369, QN => n3228);
   KEY_EXPAN0_reg_39_2_inst : FD1 port map( D => n4772, CP => CLK_I, Q => 
                           n_2370, QN => n3215);
   KEY_EXPAN0_reg_38_2_inst : FD1 port map( D => n4771, CP => CLK_I, Q => 
                           n_2371, QN => n3214);
   KEY_EXPAN0_reg_37_2_inst : FD1 port map( D => n4770, CP => CLK_I, Q => 
                           n_2372, QN => n3217);
   KEY_EXPAN0_reg_36_2_inst : FD1 port map( D => n4769, CP => CLK_I, Q => 
                           n_2373, QN => n3216);
   KEY_EXPAN0_reg_35_2_inst : FD1 port map( D => n4768, CP => CLK_I, Q => 
                           n_2374, QN => n3219);
   KEY_EXPAN0_reg_34_2_inst : FD1 port map( D => n4767, CP => CLK_I, Q => 
                           n_2375, QN => n3218);
   KEY_EXPAN0_reg_33_2_inst : FD1 port map( D => n4766, CP => CLK_I, Q => 
                           n_2376, QN => n3221);
   KEY_EXPAN0_reg_32_2_inst : FD1 port map( D => n4765, CP => CLK_I, Q => 
                           n_2377, QN => n3220);
   KEY_EXPAN0_reg_31_2_inst : FD1 port map( D => n4764, CP => CLK_I, Q => 
                           n_2378, QN => n3271);
   KEY_EXPAN0_reg_30_2_inst : FD1 port map( D => n4763, CP => CLK_I, Q => 
                           n_2379, QN => n3270);
   KEY_EXPAN0_reg_29_2_inst : FD1 port map( D => n4762, CP => CLK_I, Q => 
                           n_2380, QN => n3273);
   KEY_EXPAN0_reg_28_2_inst : FD1 port map( D => n4761, CP => CLK_I, Q => 
                           n_2381, QN => n3272);
   KEY_EXPAN0_reg_27_2_inst : FD1 port map( D => n4760, CP => CLK_I, Q => 
                           n_2382, QN => n3275);
   KEY_EXPAN0_reg_26_2_inst : FD1 port map( D => n4759, CP => CLK_I, Q => 
                           n_2383, QN => n3274);
   KEY_EXPAN0_reg_25_2_inst : FD1 port map( D => n4758, CP => CLK_I, Q => 
                           n_2384, QN => n3277);
   KEY_EXPAN0_reg_24_2_inst : FD1 port map( D => n4757, CP => CLK_I, Q => 
                           n_2385, QN => n3276);
   KEY_EXPAN0_reg_23_2_inst : FD1 port map( D => n4756, CP => CLK_I, Q => 
                           n_2386, QN => n3263);
   KEY_EXPAN0_reg_22_2_inst : FD1 port map( D => n4755, CP => CLK_I, Q => 
                           n_2387, QN => n3262);
   KEY_EXPAN0_reg_21_2_inst : FD1 port map( D => n4754, CP => CLK_I, Q => 
                           n_2388, QN => n3265);
   KEY_EXPAN0_reg_20_2_inst : FD1 port map( D => n4753, CP => CLK_I, Q => 
                           n_2389, QN => n3264);
   KEY_EXPAN0_reg_19_2_inst : FD1 port map( D => n4752, CP => CLK_I, Q => 
                           n_2390, QN => n3267);
   KEY_EXPAN0_reg_18_2_inst : FD1 port map( D => n4751, CP => CLK_I, Q => 
                           n_2391, QN => n3266);
   KEY_EXPAN0_reg_17_2_inst : FD1 port map( D => n4750, CP => CLK_I, Q => 
                           n_2392, QN => n3269);
   KEY_EXPAN0_reg_16_2_inst : FD1 port map( D => n4749, CP => CLK_I, Q => 
                           n_2393, QN => n3268);
   KEY_EXPAN0_reg_15_2_inst : FD1 port map( D => n4748, CP => CLK_I, Q => 
                           n_2394, QN => n3255);
   KEY_EXPAN0_reg_14_2_inst : FD1 port map( D => n4747, CP => CLK_I, Q => 
                           n_2395, QN => n3254);
   KEY_EXPAN0_reg_13_2_inst : FD1 port map( D => n4746, CP => CLK_I, Q => 
                           n_2396, QN => n3257);
   KEY_EXPAN0_reg_12_2_inst : FD1 port map( D => n4745, CP => CLK_I, Q => 
                           n_2397, QN => n3256);
   KEY_EXPAN0_reg_11_2_inst : FD1 port map( D => n4744, CP => CLK_I, Q => 
                           n_2398, QN => n3259);
   KEY_EXPAN0_reg_10_2_inst : FD1 port map( D => n4743, CP => CLK_I, Q => 
                           n_2399, QN => n3258);
   KEY_EXPAN0_reg_9_2_inst : FD1 port map( D => n4742, CP => CLK_I, Q => n_2400
                           , QN => n3261);
   KEY_EXPAN0_reg_8_2_inst : FD1 port map( D => n4741, CP => CLK_I, Q => n_2401
                           , QN => n3260);
   KEY_EXPAN0_reg_7_2_inst : FD1 port map( D => n4740, CP => CLK_I, Q => n_2402
                           , QN => n3247);
   KEY_EXPAN0_reg_6_2_inst : FD1 port map( D => n4739, CP => CLK_I, Q => n_2403
                           , QN => n3246);
   KEY_EXPAN0_reg_5_2_inst : FD1 port map( D => n4738, CP => CLK_I, Q => n_2404
                           , QN => n3249);
   KEY_EXPAN0_reg_4_2_inst : FD1 port map( D => n4737, CP => CLK_I, Q => n_2405
                           , QN => n3248);
   KEY_EXPAN0_reg_3_2_inst : FD1 port map( D => n4736, CP => CLK_I, Q => n_2406
                           , QN => n3251);
   KEY_EXPAN0_reg_2_2_inst : FD1 port map( D => n4735, CP => CLK_I, Q => n_2407
                           , QN => n3250);
   KEY_EXPAN0_reg_1_2_inst : FD1 port map( D => n4734, CP => CLK_I, Q => n_2408
                           , QN => n3253);
   KEY_EXPAN0_reg_0_2_inst : FD1 port map( D => n4733, CP => CLK_I, Q => n_2409
                           , QN => n3252);
   v_KEY_COL_OUT0_reg_2_inst : FD1 port map( D => n4575, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_2_port, QN => n1968);
   v_TEMP_VECTOR_reg_26_inst : FD1 port map( D => n6683, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_26_port, QN => n_2410);
   KEY_EXPAN0_reg_63_26_inst : FD1 port map( D => n6332, CP => CLK_I, Q => 
                           n_2411, QN => n3175);
   KEY_EXPAN0_reg_62_26_inst : FD1 port map( D => n6331, CP => CLK_I, Q => 
                           n_2412, QN => n3174);
   KEY_EXPAN0_reg_61_26_inst : FD1 port map( D => n6330, CP => CLK_I, Q => 
                           n_2413, QN => n3177);
   KEY_EXPAN0_reg_60_26_inst : FD1 port map( D => n6329, CP => CLK_I, Q => 
                           n_2414, QN => n3176);
   KEY_EXPAN0_reg_59_26_inst : FD1 port map( D => n6328, CP => CLK_I, Q => 
                           n_2415, QN => n3179);
   KEY_EXPAN0_reg_58_26_inst : FD1 port map( D => n6327, CP => CLK_I, Q => 
                           n_2416, QN => n3178);
   KEY_EXPAN0_reg_57_26_inst : FD1 port map( D => n6326, CP => CLK_I, Q => 
                           n_2417, QN => n3181);
   KEY_EXPAN0_reg_56_26_inst : FD1 port map( D => n6325, CP => CLK_I, Q => 
                           n_2418, QN => n3180);
   KEY_EXPAN0_reg_55_26_inst : FD1 port map( D => n6324, CP => CLK_I, Q => 
                           n_2419, QN => n3167);
   KEY_EXPAN0_reg_54_26_inst : FD1 port map( D => n6323, CP => CLK_I, Q => 
                           n_2420, QN => n3166);
   KEY_EXPAN0_reg_53_26_inst : FD1 port map( D => n6322, CP => CLK_I, Q => 
                           n_2421, QN => n3169);
   KEY_EXPAN0_reg_52_26_inst : FD1 port map( D => n6321, CP => CLK_I, Q => 
                           n_2422, QN => n3168);
   KEY_EXPAN0_reg_51_26_inst : FD1 port map( D => n6320, CP => CLK_I, Q => 
                           n_2423, QN => n3171);
   KEY_EXPAN0_reg_50_26_inst : FD1 port map( D => n6319, CP => CLK_I, Q => 
                           n_2424, QN => n3170);
   KEY_EXPAN0_reg_49_26_inst : FD1 port map( D => n6318, CP => CLK_I, Q => 
                           n_2425, QN => n3173);
   KEY_EXPAN0_reg_48_26_inst : FD1 port map( D => n6317, CP => CLK_I, Q => 
                           n_2426, QN => n3172);
   KEY_EXPAN0_reg_47_26_inst : FD1 port map( D => n6316, CP => CLK_I, Q => 
                           n_2427, QN => n3159);
   KEY_EXPAN0_reg_46_26_inst : FD1 port map( D => n6315, CP => CLK_I, Q => 
                           n_2428, QN => n3158);
   KEY_EXPAN0_reg_45_26_inst : FD1 port map( D => n6314, CP => CLK_I, Q => 
                           n_2429, QN => n3161);
   KEY_EXPAN0_reg_44_26_inst : FD1 port map( D => n6313, CP => CLK_I, Q => 
                           n_2430, QN => n3160);
   KEY_EXPAN0_reg_43_26_inst : FD1 port map( D => n6312, CP => CLK_I, Q => 
                           n_2431, QN => n3163);
   KEY_EXPAN0_reg_42_26_inst : FD1 port map( D => n6311, CP => CLK_I, Q => 
                           n_2432, QN => n3162);
   KEY_EXPAN0_reg_41_26_inst : FD1 port map( D => n6310, CP => CLK_I, Q => 
                           n_2433, QN => n3165);
   KEY_EXPAN0_reg_40_26_inst : FD1 port map( D => n6309, CP => CLK_I, Q => 
                           n_2434, QN => n3164);
   KEY_EXPAN0_reg_39_26_inst : FD1 port map( D => n6308, CP => CLK_I, Q => 
                           n_2435, QN => n3151);
   KEY_EXPAN0_reg_38_26_inst : FD1 port map( D => n6307, CP => CLK_I, Q => 
                           n_2436, QN => n3150);
   KEY_EXPAN0_reg_37_26_inst : FD1 port map( D => n6306, CP => CLK_I, Q => 
                           n_2437, QN => n3153);
   KEY_EXPAN0_reg_36_26_inst : FD1 port map( D => n6305, CP => CLK_I, Q => 
                           n_2438, QN => n3152);
   KEY_EXPAN0_reg_35_26_inst : FD1 port map( D => n6304, CP => CLK_I, Q => 
                           n_2439, QN => n3155);
   KEY_EXPAN0_reg_34_26_inst : FD1 port map( D => n6303, CP => CLK_I, Q => 
                           n_2440, QN => n3154);
   KEY_EXPAN0_reg_33_26_inst : FD1 port map( D => n6302, CP => CLK_I, Q => 
                           n_2441, QN => n3157);
   KEY_EXPAN0_reg_32_26_inst : FD1 port map( D => n6301, CP => CLK_I, Q => 
                           n_2442, QN => n3156);
   KEY_EXPAN0_reg_31_26_inst : FD1 port map( D => n6300, CP => CLK_I, Q => 
                           n_2443, QN => n3207);
   KEY_EXPAN0_reg_30_26_inst : FD1 port map( D => n6299, CP => CLK_I, Q => 
                           n_2444, QN => n3206);
   KEY_EXPAN0_reg_29_26_inst : FD1 port map( D => n6298, CP => CLK_I, Q => 
                           n_2445, QN => n3209);
   KEY_EXPAN0_reg_28_26_inst : FD1 port map( D => n6297, CP => CLK_I, Q => 
                           n_2446, QN => n3208);
   KEY_EXPAN0_reg_27_26_inst : FD1 port map( D => n6296, CP => CLK_I, Q => 
                           n_2447, QN => n3211);
   KEY_EXPAN0_reg_26_26_inst : FD1 port map( D => n6295, CP => CLK_I, Q => 
                           n_2448, QN => n3210);
   KEY_EXPAN0_reg_25_26_inst : FD1 port map( D => n6294, CP => CLK_I, Q => 
                           n_2449, QN => n3213);
   KEY_EXPAN0_reg_24_26_inst : FD1 port map( D => n6293, CP => CLK_I, Q => 
                           n_2450, QN => n3212);
   KEY_EXPAN0_reg_23_26_inst : FD1 port map( D => n6292, CP => CLK_I, Q => 
                           n_2451, QN => n3199);
   KEY_EXPAN0_reg_22_26_inst : FD1 port map( D => n6291, CP => CLK_I, Q => 
                           n_2452, QN => n3198);
   KEY_EXPAN0_reg_21_26_inst : FD1 port map( D => n6290, CP => CLK_I, Q => 
                           n_2453, QN => n3201);
   KEY_EXPAN0_reg_20_26_inst : FD1 port map( D => n6289, CP => CLK_I, Q => 
                           n_2454, QN => n3200);
   KEY_EXPAN0_reg_19_26_inst : FD1 port map( D => n6288, CP => CLK_I, Q => 
                           n_2455, QN => n3203);
   KEY_EXPAN0_reg_18_26_inst : FD1 port map( D => n6287, CP => CLK_I, Q => 
                           n_2456, QN => n3202);
   KEY_EXPAN0_reg_17_26_inst : FD1 port map( D => n6286, CP => CLK_I, Q => 
                           n_2457, QN => n3205);
   KEY_EXPAN0_reg_16_26_inst : FD1 port map( D => n6285, CP => CLK_I, Q => 
                           n_2458, QN => n3204);
   KEY_EXPAN0_reg_15_26_inst : FD1 port map( D => n6284, CP => CLK_I, Q => 
                           n_2459, QN => n3191);
   KEY_EXPAN0_reg_14_26_inst : FD1 port map( D => n6283, CP => CLK_I, Q => 
                           n_2460, QN => n3190);
   KEY_EXPAN0_reg_13_26_inst : FD1 port map( D => n6282, CP => CLK_I, Q => 
                           n_2461, QN => n3193);
   KEY_EXPAN0_reg_12_26_inst : FD1 port map( D => n6281, CP => CLK_I, Q => 
                           n_2462, QN => n3192);
   KEY_EXPAN0_reg_11_26_inst : FD1 port map( D => n6280, CP => CLK_I, Q => 
                           n_2463, QN => n3195);
   KEY_EXPAN0_reg_10_26_inst : FD1 port map( D => n6279, CP => CLK_I, Q => 
                           n_2464, QN => n3194);
   KEY_EXPAN0_reg_9_26_inst : FD1 port map( D => n6278, CP => CLK_I, Q => 
                           n_2465, QN => n3197);
   KEY_EXPAN0_reg_8_26_inst : FD1 port map( D => n6277, CP => CLK_I, Q => 
                           n_2466, QN => n3196);
   KEY_EXPAN0_reg_7_26_inst : FD1 port map( D => n6276, CP => CLK_I, Q => 
                           n_2467, QN => n3183);
   KEY_EXPAN0_reg_6_26_inst : FD1 port map( D => n6275, CP => CLK_I, Q => 
                           n_2468, QN => n3182);
   KEY_EXPAN0_reg_5_26_inst : FD1 port map( D => n6274, CP => CLK_I, Q => 
                           n_2469, QN => n3185);
   KEY_EXPAN0_reg_4_26_inst : FD1 port map( D => n6273, CP => CLK_I, Q => 
                           n_2470, QN => n3184);
   KEY_EXPAN0_reg_3_26_inst : FD1 port map( D => n6272, CP => CLK_I, Q => 
                           n_2471, QN => n3187);
   KEY_EXPAN0_reg_2_26_inst : FD1 port map( D => n6271, CP => CLK_I, Q => 
                           n_2472, QN => n3186);
   KEY_EXPAN0_reg_1_26_inst : FD1 port map( D => n6270, CP => CLK_I, Q => 
                           n_2473, QN => n3189);
   KEY_EXPAN0_reg_0_26_inst : FD1 port map( D => n6269, CP => CLK_I, Q => 
                           n_2474, QN => n3188);
   v_KEY_COL_OUT0_reg_26_inst : FD1 port map( D => n4574, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_26_port, QN => n1999);
   v_TEMP_VECTOR_reg_18_inst : FD1 port map( D => n6691, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_18_port, QN => n_2475);
   KEY_EXPAN0_reg_63_18_inst : FD1 port map( D => n5820, CP => CLK_I, Q => 
                           n_2476, QN => n3111);
   KEY_EXPAN0_reg_62_18_inst : FD1 port map( D => n5819, CP => CLK_I, Q => 
                           n_2477, QN => n3110);
   KEY_EXPAN0_reg_61_18_inst : FD1 port map( D => n5818, CP => CLK_I, Q => 
                           n_2478, QN => n3113);
   KEY_EXPAN0_reg_60_18_inst : FD1 port map( D => n5817, CP => CLK_I, Q => 
                           n_2479, QN => n3112);
   KEY_EXPAN0_reg_59_18_inst : FD1 port map( D => n5816, CP => CLK_I, Q => 
                           n_2480, QN => n3115);
   KEY_EXPAN0_reg_58_18_inst : FD1 port map( D => n5815, CP => CLK_I, Q => 
                           n_2481, QN => n3114);
   KEY_EXPAN0_reg_57_18_inst : FD1 port map( D => n5814, CP => CLK_I, Q => 
                           n_2482, QN => n3117);
   KEY_EXPAN0_reg_56_18_inst : FD1 port map( D => n5813, CP => CLK_I, Q => 
                           n_2483, QN => n3116);
   KEY_EXPAN0_reg_55_18_inst : FD1 port map( D => n5812, CP => CLK_I, Q => 
                           n_2484, QN => n3103);
   KEY_EXPAN0_reg_54_18_inst : FD1 port map( D => n5811, CP => CLK_I, Q => 
                           n_2485, QN => n3102);
   KEY_EXPAN0_reg_53_18_inst : FD1 port map( D => n5810, CP => CLK_I, Q => 
                           n_2486, QN => n3105);
   KEY_EXPAN0_reg_52_18_inst : FD1 port map( D => n5809, CP => CLK_I, Q => 
                           n_2487, QN => n3104);
   KEY_EXPAN0_reg_51_18_inst : FD1 port map( D => n5808, CP => CLK_I, Q => 
                           n_2488, QN => n3107);
   KEY_EXPAN0_reg_50_18_inst : FD1 port map( D => n5807, CP => CLK_I, Q => 
                           n_2489, QN => n3106);
   KEY_EXPAN0_reg_49_18_inst : FD1 port map( D => n5806, CP => CLK_I, Q => 
                           n_2490, QN => n3109);
   KEY_EXPAN0_reg_48_18_inst : FD1 port map( D => n5805, CP => CLK_I, Q => 
                           n_2491, QN => n3108);
   KEY_EXPAN0_reg_47_18_inst : FD1 port map( D => n5804, CP => CLK_I, Q => 
                           n_2492, QN => n3095);
   KEY_EXPAN0_reg_46_18_inst : FD1 port map( D => n5803, CP => CLK_I, Q => 
                           n_2493, QN => n3094);
   KEY_EXPAN0_reg_45_18_inst : FD1 port map( D => n5802, CP => CLK_I, Q => 
                           n_2494, QN => n3097);
   KEY_EXPAN0_reg_44_18_inst : FD1 port map( D => n5801, CP => CLK_I, Q => 
                           n_2495, QN => n3096);
   KEY_EXPAN0_reg_43_18_inst : FD1 port map( D => n5800, CP => CLK_I, Q => 
                           n_2496, QN => n3099);
   KEY_EXPAN0_reg_42_18_inst : FD1 port map( D => n5799, CP => CLK_I, Q => 
                           n_2497, QN => n3098);
   KEY_EXPAN0_reg_41_18_inst : FD1 port map( D => n5798, CP => CLK_I, Q => 
                           n_2498, QN => n3101);
   KEY_EXPAN0_reg_40_18_inst : FD1 port map( D => n5797, CP => CLK_I, Q => 
                           n_2499, QN => n3100);
   KEY_EXPAN0_reg_39_18_inst : FD1 port map( D => n5796, CP => CLK_I, Q => 
                           n_2500, QN => n3087);
   KEY_EXPAN0_reg_38_18_inst : FD1 port map( D => n5795, CP => CLK_I, Q => 
                           n_2501, QN => n3086);
   KEY_EXPAN0_reg_37_18_inst : FD1 port map( D => n5794, CP => CLK_I, Q => 
                           n_2502, QN => n3089);
   KEY_EXPAN0_reg_36_18_inst : FD1 port map( D => n5793, CP => CLK_I, Q => 
                           n_2503, QN => n3088);
   KEY_EXPAN0_reg_35_18_inst : FD1 port map( D => n5792, CP => CLK_I, Q => 
                           n_2504, QN => n3091);
   KEY_EXPAN0_reg_34_18_inst : FD1 port map( D => n5791, CP => CLK_I, Q => 
                           n_2505, QN => n3090);
   KEY_EXPAN0_reg_33_18_inst : FD1 port map( D => n5790, CP => CLK_I, Q => 
                           n_2506, QN => n3093);
   KEY_EXPAN0_reg_32_18_inst : FD1 port map( D => n5789, CP => CLK_I, Q => 
                           n_2507, QN => n3092);
   KEY_EXPAN0_reg_31_18_inst : FD1 port map( D => n5788, CP => CLK_I, Q => 
                           n_2508, QN => n3143);
   KEY_EXPAN0_reg_30_18_inst : FD1 port map( D => n5787, CP => CLK_I, Q => 
                           n_2509, QN => n3142);
   KEY_EXPAN0_reg_29_18_inst : FD1 port map( D => n5786, CP => CLK_I, Q => 
                           n_2510, QN => n3145);
   KEY_EXPAN0_reg_28_18_inst : FD1 port map( D => n5785, CP => CLK_I, Q => 
                           n_2511, QN => n3144);
   KEY_EXPAN0_reg_27_18_inst : FD1 port map( D => n5784, CP => CLK_I, Q => 
                           n_2512, QN => n3147);
   KEY_EXPAN0_reg_26_18_inst : FD1 port map( D => n5783, CP => CLK_I, Q => 
                           n_2513, QN => n3146);
   KEY_EXPAN0_reg_25_18_inst : FD1 port map( D => n5782, CP => CLK_I, Q => 
                           n_2514, QN => n3149);
   KEY_EXPAN0_reg_24_18_inst : FD1 port map( D => n5781, CP => CLK_I, Q => 
                           n_2515, QN => n3148);
   KEY_EXPAN0_reg_23_18_inst : FD1 port map( D => n5780, CP => CLK_I, Q => 
                           n_2516, QN => n3135);
   KEY_EXPAN0_reg_22_18_inst : FD1 port map( D => n5779, CP => CLK_I, Q => 
                           n_2517, QN => n3134);
   KEY_EXPAN0_reg_21_18_inst : FD1 port map( D => n5778, CP => CLK_I, Q => 
                           n_2518, QN => n3137);
   KEY_EXPAN0_reg_20_18_inst : FD1 port map( D => n5777, CP => CLK_I, Q => 
                           n_2519, QN => n3136);
   KEY_EXPAN0_reg_19_18_inst : FD1 port map( D => n5776, CP => CLK_I, Q => 
                           n_2520, QN => n3139);
   KEY_EXPAN0_reg_18_18_inst : FD1 port map( D => n5775, CP => CLK_I, Q => 
                           n_2521, QN => n3138);
   KEY_EXPAN0_reg_17_18_inst : FD1 port map( D => n5774, CP => CLK_I, Q => 
                           n_2522, QN => n3141);
   KEY_EXPAN0_reg_16_18_inst : FD1 port map( D => n5773, CP => CLK_I, Q => 
                           n_2523, QN => n3140);
   KEY_EXPAN0_reg_15_18_inst : FD1 port map( D => n5772, CP => CLK_I, Q => 
                           n_2524, QN => n3127);
   KEY_EXPAN0_reg_14_18_inst : FD1 port map( D => n5771, CP => CLK_I, Q => 
                           n_2525, QN => n3126);
   KEY_EXPAN0_reg_13_18_inst : FD1 port map( D => n5770, CP => CLK_I, Q => 
                           n_2526, QN => n3129);
   KEY_EXPAN0_reg_12_18_inst : FD1 port map( D => n5769, CP => CLK_I, Q => 
                           n_2527, QN => n3128);
   KEY_EXPAN0_reg_11_18_inst : FD1 port map( D => n5768, CP => CLK_I, Q => 
                           n_2528, QN => n3131);
   KEY_EXPAN0_reg_10_18_inst : FD1 port map( D => n5767, CP => CLK_I, Q => 
                           n_2529, QN => n3130);
   KEY_EXPAN0_reg_9_18_inst : FD1 port map( D => n5766, CP => CLK_I, Q => 
                           n_2530, QN => n3133);
   KEY_EXPAN0_reg_8_18_inst : FD1 port map( D => n5765, CP => CLK_I, Q => 
                           n_2531, QN => n3132);
   KEY_EXPAN0_reg_7_18_inst : FD1 port map( D => n5764, CP => CLK_I, Q => 
                           n_2532, QN => n3119);
   KEY_EXPAN0_reg_6_18_inst : FD1 port map( D => n5763, CP => CLK_I, Q => 
                           n_2533, QN => n3118);
   KEY_EXPAN0_reg_5_18_inst : FD1 port map( D => n5762, CP => CLK_I, Q => 
                           n_2534, QN => n3121);
   KEY_EXPAN0_reg_4_18_inst : FD1 port map( D => n5761, CP => CLK_I, Q => 
                           n_2535, QN => n3120);
   KEY_EXPAN0_reg_3_18_inst : FD1 port map( D => n5760, CP => CLK_I, Q => 
                           n_2536, QN => n3123);
   KEY_EXPAN0_reg_2_18_inst : FD1 port map( D => n5759, CP => CLK_I, Q => 
                           n_2537, QN => n3122);
   KEY_EXPAN0_reg_1_18_inst : FD1 port map( D => n5758, CP => CLK_I, Q => 
                           n_2538, QN => n3125);
   KEY_EXPAN0_reg_0_18_inst : FD1 port map( D => n5757, CP => CLK_I, Q => 
                           n_2539, QN => n3124);
   v_KEY_COL_OUT0_reg_18_inst : FD1 port map( D => n4573, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_18_port, QN => n1956);
   v_TEMP_VECTOR_reg_10_inst : FD1 port map( D => n6699, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_10_port, QN => n_2540);
   KEY_EXPAN0_reg_63_10_inst : FD1 port map( D => n5308, CP => CLK_I, Q => 
                           n_2541, QN => n3047);
   KEY_EXPAN0_reg_62_10_inst : FD1 port map( D => n5307, CP => CLK_I, Q => 
                           n_2542, QN => n3046);
   KEY_EXPAN0_reg_61_10_inst : FD1 port map( D => n5306, CP => CLK_I, Q => 
                           n_2543, QN => n3049);
   KEY_EXPAN0_reg_60_10_inst : FD1 port map( D => n5305, CP => CLK_I, Q => 
                           n_2544, QN => n3048);
   KEY_EXPAN0_reg_59_10_inst : FD1 port map( D => n5304, CP => CLK_I, Q => 
                           n_2545, QN => n3051);
   KEY_EXPAN0_reg_58_10_inst : FD1 port map( D => n5303, CP => CLK_I, Q => 
                           n_2546, QN => n3050);
   KEY_EXPAN0_reg_57_10_inst : FD1 port map( D => n5302, CP => CLK_I, Q => 
                           n_2547, QN => n3053);
   KEY_EXPAN0_reg_56_10_inst : FD1 port map( D => n5301, CP => CLK_I, Q => 
                           n_2548, QN => n3052);
   KEY_EXPAN0_reg_55_10_inst : FD1 port map( D => n5300, CP => CLK_I, Q => 
                           n_2549, QN => n3039);
   KEY_EXPAN0_reg_54_10_inst : FD1 port map( D => n5299, CP => CLK_I, Q => 
                           n_2550, QN => n3038);
   KEY_EXPAN0_reg_53_10_inst : FD1 port map( D => n5298, CP => CLK_I, Q => 
                           n_2551, QN => n3041);
   KEY_EXPAN0_reg_52_10_inst : FD1 port map( D => n5297, CP => CLK_I, Q => 
                           n_2552, QN => n3040);
   KEY_EXPAN0_reg_51_10_inst : FD1 port map( D => n5296, CP => CLK_I, Q => 
                           n_2553, QN => n3043);
   KEY_EXPAN0_reg_50_10_inst : FD1 port map( D => n5295, CP => CLK_I, Q => 
                           n_2554, QN => n3042);
   KEY_EXPAN0_reg_49_10_inst : FD1 port map( D => n5294, CP => CLK_I, Q => 
                           n_2555, QN => n3045);
   KEY_EXPAN0_reg_48_10_inst : FD1 port map( D => n5293, CP => CLK_I, Q => 
                           n_2556, QN => n3044);
   KEY_EXPAN0_reg_47_10_inst : FD1 port map( D => n5292, CP => CLK_I, Q => 
                           n_2557, QN => n3031);
   KEY_EXPAN0_reg_46_10_inst : FD1 port map( D => n5291, CP => CLK_I, Q => 
                           n_2558, QN => n3030);
   KEY_EXPAN0_reg_45_10_inst : FD1 port map( D => n5290, CP => CLK_I, Q => 
                           n_2559, QN => n3033);
   KEY_EXPAN0_reg_44_10_inst : FD1 port map( D => n5289, CP => CLK_I, Q => 
                           n_2560, QN => n3032);
   KEY_EXPAN0_reg_43_10_inst : FD1 port map( D => n5288, CP => CLK_I, Q => 
                           n_2561, QN => n3035);
   KEY_EXPAN0_reg_42_10_inst : FD1 port map( D => n5287, CP => CLK_I, Q => 
                           n_2562, QN => n3034);
   KEY_EXPAN0_reg_41_10_inst : FD1 port map( D => n5286, CP => CLK_I, Q => 
                           n_2563, QN => n3037);
   KEY_EXPAN0_reg_40_10_inst : FD1 port map( D => n5285, CP => CLK_I, Q => 
                           n_2564, QN => n3036);
   KEY_EXPAN0_reg_39_10_inst : FD1 port map( D => n5284, CP => CLK_I, Q => 
                           n_2565, QN => n3023);
   KEY_EXPAN0_reg_38_10_inst : FD1 port map( D => n5283, CP => CLK_I, Q => 
                           n_2566, QN => n3022);
   KEY_EXPAN0_reg_37_10_inst : FD1 port map( D => n5282, CP => CLK_I, Q => 
                           n_2567, QN => n3025);
   KEY_EXPAN0_reg_36_10_inst : FD1 port map( D => n5281, CP => CLK_I, Q => 
                           n_2568, QN => n3024);
   KEY_EXPAN0_reg_35_10_inst : FD1 port map( D => n5280, CP => CLK_I, Q => 
                           n_2569, QN => n3027);
   KEY_EXPAN0_reg_34_10_inst : FD1 port map( D => n5279, CP => CLK_I, Q => 
                           n_2570, QN => n3026);
   KEY_EXPAN0_reg_33_10_inst : FD1 port map( D => n5278, CP => CLK_I, Q => 
                           n_2571, QN => n3029);
   KEY_EXPAN0_reg_32_10_inst : FD1 port map( D => n5277, CP => CLK_I, Q => 
                           n_2572, QN => n3028);
   KEY_EXPAN0_reg_31_10_inst : FD1 port map( D => n5276, CP => CLK_I, Q => 
                           n_2573, QN => n3079);
   KEY_EXPAN0_reg_30_10_inst : FD1 port map( D => n5275, CP => CLK_I, Q => 
                           n_2574, QN => n3078);
   KEY_EXPAN0_reg_29_10_inst : FD1 port map( D => n5274, CP => CLK_I, Q => 
                           n_2575, QN => n3081);
   KEY_EXPAN0_reg_28_10_inst : FD1 port map( D => n5273, CP => CLK_I, Q => 
                           n_2576, QN => n3080);
   KEY_EXPAN0_reg_27_10_inst : FD1 port map( D => n5272, CP => CLK_I, Q => 
                           n_2577, QN => n3083);
   KEY_EXPAN0_reg_26_10_inst : FD1 port map( D => n5271, CP => CLK_I, Q => 
                           n_2578, QN => n3082);
   KEY_EXPAN0_reg_25_10_inst : FD1 port map( D => n5270, CP => CLK_I, Q => 
                           n_2579, QN => n3085);
   KEY_EXPAN0_reg_24_10_inst : FD1 port map( D => n5269, CP => CLK_I, Q => 
                           n_2580, QN => n3084);
   KEY_EXPAN0_reg_23_10_inst : FD1 port map( D => n5268, CP => CLK_I, Q => 
                           n_2581, QN => n3071);
   KEY_EXPAN0_reg_22_10_inst : FD1 port map( D => n5267, CP => CLK_I, Q => 
                           n_2582, QN => n3070);
   KEY_EXPAN0_reg_21_10_inst : FD1 port map( D => n5266, CP => CLK_I, Q => 
                           n_2583, QN => n3073);
   KEY_EXPAN0_reg_20_10_inst : FD1 port map( D => n5265, CP => CLK_I, Q => 
                           n_2584, QN => n3072);
   KEY_EXPAN0_reg_19_10_inst : FD1 port map( D => n5264, CP => CLK_I, Q => 
                           n_2585, QN => n3075);
   KEY_EXPAN0_reg_18_10_inst : FD1 port map( D => n5263, CP => CLK_I, Q => 
                           n_2586, QN => n3074);
   KEY_EXPAN0_reg_17_10_inst : FD1 port map( D => n5262, CP => CLK_I, Q => 
                           n_2587, QN => n3077);
   KEY_EXPAN0_reg_16_10_inst : FD1 port map( D => n5261, CP => CLK_I, Q => 
                           n_2588, QN => n3076);
   KEY_EXPAN0_reg_15_10_inst : FD1 port map( D => n5260, CP => CLK_I, Q => 
                           n_2589, QN => n3063);
   KEY_EXPAN0_reg_14_10_inst : FD1 port map( D => n5259, CP => CLK_I, Q => 
                           n_2590, QN => n3062);
   KEY_EXPAN0_reg_13_10_inst : FD1 port map( D => n5258, CP => CLK_I, Q => 
                           n_2591, QN => n3065);
   KEY_EXPAN0_reg_12_10_inst : FD1 port map( D => n5257, CP => CLK_I, Q => 
                           n_2592, QN => n3064);
   KEY_EXPAN0_reg_11_10_inst : FD1 port map( D => n5256, CP => CLK_I, Q => 
                           n_2593, QN => n3067);
   KEY_EXPAN0_reg_10_10_inst : FD1 port map( D => n5255, CP => CLK_I, Q => 
                           n_2594, QN => n3066);
   KEY_EXPAN0_reg_9_10_inst : FD1 port map( D => n5254, CP => CLK_I, Q => 
                           n_2595, QN => n3069);
   KEY_EXPAN0_reg_8_10_inst : FD1 port map( D => n5253, CP => CLK_I, Q => 
                           n_2596, QN => n3068);
   KEY_EXPAN0_reg_7_10_inst : FD1 port map( D => n5252, CP => CLK_I, Q => 
                           n_2597, QN => n3055);
   KEY_EXPAN0_reg_6_10_inst : FD1 port map( D => n5251, CP => CLK_I, Q => 
                           n_2598, QN => n3054);
   KEY_EXPAN0_reg_5_10_inst : FD1 port map( D => n5250, CP => CLK_I, Q => 
                           n_2599, QN => n3057);
   KEY_EXPAN0_reg_4_10_inst : FD1 port map( D => n5249, CP => CLK_I, Q => 
                           n_2600, QN => n3056);
   KEY_EXPAN0_reg_3_10_inst : FD1 port map( D => n5248, CP => CLK_I, Q => 
                           n_2601, QN => n3059);
   KEY_EXPAN0_reg_2_10_inst : FD1 port map( D => n5247, CP => CLK_I, Q => 
                           n_2602, QN => n3058);
   KEY_EXPAN0_reg_1_10_inst : FD1 port map( D => n5246, CP => CLK_I, Q => 
                           n_2603, QN => n3061);
   KEY_EXPAN0_reg_0_10_inst : FD1 port map( D => n5245, CP => CLK_I, Q => 
                           n_2604, QN => n3060);
   v_KEY_COL_OUT0_reg_10_inst : FD1 port map( D => n4572, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_10_port, QN => n1922);
   v_TEMP_VECTOR_reg_1_inst : FD1 port map( D => n6708, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_1_port, QN => n_2605);
   KEY_EXPAN0_reg_63_1_inst : FD1 port map( D => n4732, CP => CLK_I, Q => 
                           n_2606, QN => n2983);
   KEY_EXPAN0_reg_62_1_inst : FD1 port map( D => n4731, CP => CLK_I, Q => 
                           n_2607, QN => n2982);
   KEY_EXPAN0_reg_61_1_inst : FD1 port map( D => n4730, CP => CLK_I, Q => 
                           n_2608, QN => n2985);
   KEY_EXPAN0_reg_60_1_inst : FD1 port map( D => n4729, CP => CLK_I, Q => 
                           n_2609, QN => n2984);
   KEY_EXPAN0_reg_59_1_inst : FD1 port map( D => n4728, CP => CLK_I, Q => 
                           n_2610, QN => n2987);
   KEY_EXPAN0_reg_58_1_inst : FD1 port map( D => n4727, CP => CLK_I, Q => 
                           n_2611, QN => n2986);
   KEY_EXPAN0_reg_57_1_inst : FD1 port map( D => n4726, CP => CLK_I, Q => 
                           n_2612, QN => n2989);
   KEY_EXPAN0_reg_56_1_inst : FD1 port map( D => n4725, CP => CLK_I, Q => 
                           n_2613, QN => n2988);
   KEY_EXPAN0_reg_55_1_inst : FD1 port map( D => n4724, CP => CLK_I, Q => 
                           n_2614, QN => n2975);
   KEY_EXPAN0_reg_54_1_inst : FD1 port map( D => n4723, CP => CLK_I, Q => 
                           n_2615, QN => n2974);
   KEY_EXPAN0_reg_53_1_inst : FD1 port map( D => n4722, CP => CLK_I, Q => 
                           n_2616, QN => n2977);
   KEY_EXPAN0_reg_52_1_inst : FD1 port map( D => n4721, CP => CLK_I, Q => 
                           n_2617, QN => n2976);
   KEY_EXPAN0_reg_51_1_inst : FD1 port map( D => n4720, CP => CLK_I, Q => 
                           n_2618, QN => n2979);
   KEY_EXPAN0_reg_50_1_inst : FD1 port map( D => n4719, CP => CLK_I, Q => 
                           n_2619, QN => n2978);
   KEY_EXPAN0_reg_49_1_inst : FD1 port map( D => n4718, CP => CLK_I, Q => 
                           n_2620, QN => n2981);
   KEY_EXPAN0_reg_48_1_inst : FD1 port map( D => n4717, CP => CLK_I, Q => 
                           n_2621, QN => n2980);
   KEY_EXPAN0_reg_47_1_inst : FD1 port map( D => n4716, CP => CLK_I, Q => 
                           n_2622, QN => n2967);
   KEY_EXPAN0_reg_46_1_inst : FD1 port map( D => n4715, CP => CLK_I, Q => 
                           n_2623, QN => n2966);
   KEY_EXPAN0_reg_45_1_inst : FD1 port map( D => n4714, CP => CLK_I, Q => 
                           n_2624, QN => n2969);
   KEY_EXPAN0_reg_44_1_inst : FD1 port map( D => n4713, CP => CLK_I, Q => 
                           n_2625, QN => n2968);
   KEY_EXPAN0_reg_43_1_inst : FD1 port map( D => n4712, CP => CLK_I, Q => 
                           n_2626, QN => n2971);
   KEY_EXPAN0_reg_42_1_inst : FD1 port map( D => n4711, CP => CLK_I, Q => 
                           n_2627, QN => n2970);
   KEY_EXPAN0_reg_41_1_inst : FD1 port map( D => n4710, CP => CLK_I, Q => 
                           n_2628, QN => n2973);
   KEY_EXPAN0_reg_40_1_inst : FD1 port map( D => n4709, CP => CLK_I, Q => 
                           n_2629, QN => n2972);
   KEY_EXPAN0_reg_39_1_inst : FD1 port map( D => n4708, CP => CLK_I, Q => 
                           n_2630, QN => n2959);
   KEY_EXPAN0_reg_38_1_inst : FD1 port map( D => n4707, CP => CLK_I, Q => 
                           n_2631, QN => n2958);
   KEY_EXPAN0_reg_37_1_inst : FD1 port map( D => n4706, CP => CLK_I, Q => 
                           n_2632, QN => n2961);
   KEY_EXPAN0_reg_36_1_inst : FD1 port map( D => n4705, CP => CLK_I, Q => 
                           n_2633, QN => n2960);
   KEY_EXPAN0_reg_35_1_inst : FD1 port map( D => n4704, CP => CLK_I, Q => 
                           n_2634, QN => n2963);
   KEY_EXPAN0_reg_34_1_inst : FD1 port map( D => n4703, CP => CLK_I, Q => 
                           n_2635, QN => n2962);
   KEY_EXPAN0_reg_33_1_inst : FD1 port map( D => n4702, CP => CLK_I, Q => 
                           n_2636, QN => n2965);
   KEY_EXPAN0_reg_32_1_inst : FD1 port map( D => n4701, CP => CLK_I, Q => 
                           n_2637, QN => n2964);
   KEY_EXPAN0_reg_31_1_inst : FD1 port map( D => n4700, CP => CLK_I, Q => 
                           n_2638, QN => n3015);
   KEY_EXPAN0_reg_30_1_inst : FD1 port map( D => n4699, CP => CLK_I, Q => 
                           n_2639, QN => n3014);
   KEY_EXPAN0_reg_29_1_inst : FD1 port map( D => n4698, CP => CLK_I, Q => 
                           n_2640, QN => n3017);
   KEY_EXPAN0_reg_28_1_inst : FD1 port map( D => n4697, CP => CLK_I, Q => 
                           n_2641, QN => n3016);
   KEY_EXPAN0_reg_27_1_inst : FD1 port map( D => n4696, CP => CLK_I, Q => 
                           n_2642, QN => n3019);
   KEY_EXPAN0_reg_26_1_inst : FD1 port map( D => n4695, CP => CLK_I, Q => 
                           n_2643, QN => n3018);
   KEY_EXPAN0_reg_25_1_inst : FD1 port map( D => n4694, CP => CLK_I, Q => 
                           n_2644, QN => n3021);
   KEY_EXPAN0_reg_24_1_inst : FD1 port map( D => n4693, CP => CLK_I, Q => 
                           n_2645, QN => n3020);
   KEY_EXPAN0_reg_23_1_inst : FD1 port map( D => n4692, CP => CLK_I, Q => 
                           n_2646, QN => n3007);
   KEY_EXPAN0_reg_22_1_inst : FD1 port map( D => n4691, CP => CLK_I, Q => 
                           n_2647, QN => n3006);
   KEY_EXPAN0_reg_21_1_inst : FD1 port map( D => n4690, CP => CLK_I, Q => 
                           n_2648, QN => n3009);
   KEY_EXPAN0_reg_20_1_inst : FD1 port map( D => n4689, CP => CLK_I, Q => 
                           n_2649, QN => n3008);
   KEY_EXPAN0_reg_19_1_inst : FD1 port map( D => n4688, CP => CLK_I, Q => 
                           n_2650, QN => n3011);
   KEY_EXPAN0_reg_18_1_inst : FD1 port map( D => n4687, CP => CLK_I, Q => 
                           n_2651, QN => n3010);
   KEY_EXPAN0_reg_17_1_inst : FD1 port map( D => n4686, CP => CLK_I, Q => 
                           n_2652, QN => n3013);
   KEY_EXPAN0_reg_16_1_inst : FD1 port map( D => n4685, CP => CLK_I, Q => 
                           n_2653, QN => n3012);
   KEY_EXPAN0_reg_15_1_inst : FD1 port map( D => n4684, CP => CLK_I, Q => 
                           n_2654, QN => n2999);
   KEY_EXPAN0_reg_14_1_inst : FD1 port map( D => n4683, CP => CLK_I, Q => 
                           n_2655, QN => n2998);
   KEY_EXPAN0_reg_13_1_inst : FD1 port map( D => n4682, CP => CLK_I, Q => 
                           n_2656, QN => n3001);
   KEY_EXPAN0_reg_12_1_inst : FD1 port map( D => n4681, CP => CLK_I, Q => 
                           n_2657, QN => n3000);
   KEY_EXPAN0_reg_11_1_inst : FD1 port map( D => n4680, CP => CLK_I, Q => 
                           n_2658, QN => n3003);
   KEY_EXPAN0_reg_10_1_inst : FD1 port map( D => n4679, CP => CLK_I, Q => 
                           n_2659, QN => n3002);
   KEY_EXPAN0_reg_9_1_inst : FD1 port map( D => n4678, CP => CLK_I, Q => n_2660
                           , QN => n3005);
   KEY_EXPAN0_reg_8_1_inst : FD1 port map( D => n4677, CP => CLK_I, Q => n_2661
                           , QN => n3004);
   KEY_EXPAN0_reg_7_1_inst : FD1 port map( D => n4676, CP => CLK_I, Q => n_2662
                           , QN => n2991);
   KEY_EXPAN0_reg_6_1_inst : FD1 port map( D => n4675, CP => CLK_I, Q => n_2663
                           , QN => n2990);
   KEY_EXPAN0_reg_5_1_inst : FD1 port map( D => n4674, CP => CLK_I, Q => n_2664
                           , QN => n2993);
   KEY_EXPAN0_reg_4_1_inst : FD1 port map( D => n4673, CP => CLK_I, Q => n_2665
                           , QN => n2992);
   KEY_EXPAN0_reg_3_1_inst : FD1 port map( D => n4672, CP => CLK_I, Q => n_2666
                           , QN => n2995);
   KEY_EXPAN0_reg_2_1_inst : FD1 port map( D => n4671, CP => CLK_I, Q => n_2667
                           , QN => n2994);
   KEY_EXPAN0_reg_1_1_inst : FD1 port map( D => n4670, CP => CLK_I, Q => n_2668
                           , QN => n2997);
   KEY_EXPAN0_reg_0_1_inst : FD1 port map( D => n4669, CP => CLK_I, Q => n_2669
                           , QN => n2996);
   v_KEY_COL_OUT0_reg_1_inst : FD1 port map( D => n4571, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_1_port, QN => n1966);
   v_TEMP_VECTOR_reg_25_inst : FD1 port map( D => n6684, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_25_port, QN => n_2670);
   KEY_EXPAN0_reg_63_25_inst : FD1 port map( D => n6268, CP => CLK_I, Q => 
                           n_2671, QN => n2919);
   KEY_EXPAN0_reg_62_25_inst : FD1 port map( D => n6267, CP => CLK_I, Q => 
                           n_2672, QN => n2918);
   KEY_EXPAN0_reg_61_25_inst : FD1 port map( D => n6266, CP => CLK_I, Q => 
                           n_2673, QN => n2921);
   KEY_EXPAN0_reg_60_25_inst : FD1 port map( D => n6265, CP => CLK_I, Q => 
                           n_2674, QN => n2920);
   KEY_EXPAN0_reg_59_25_inst : FD1 port map( D => n6264, CP => CLK_I, Q => 
                           n_2675, QN => n2923);
   KEY_EXPAN0_reg_58_25_inst : FD1 port map( D => n6263, CP => CLK_I, Q => 
                           n_2676, QN => n2922);
   KEY_EXPAN0_reg_57_25_inst : FD1 port map( D => n6262, CP => CLK_I, Q => 
                           n_2677, QN => n2925);
   KEY_EXPAN0_reg_56_25_inst : FD1 port map( D => n6261, CP => CLK_I, Q => 
                           n_2678, QN => n2924);
   KEY_EXPAN0_reg_55_25_inst : FD1 port map( D => n6260, CP => CLK_I, Q => 
                           n_2679, QN => n2911);
   KEY_EXPAN0_reg_54_25_inst : FD1 port map( D => n6259, CP => CLK_I, Q => 
                           n_2680, QN => n2910);
   KEY_EXPAN0_reg_53_25_inst : FD1 port map( D => n6258, CP => CLK_I, Q => 
                           n_2681, QN => n2913);
   KEY_EXPAN0_reg_52_25_inst : FD1 port map( D => n6257, CP => CLK_I, Q => 
                           n_2682, QN => n2912);
   KEY_EXPAN0_reg_51_25_inst : FD1 port map( D => n6256, CP => CLK_I, Q => 
                           n_2683, QN => n2915);
   KEY_EXPAN0_reg_50_25_inst : FD1 port map( D => n6255, CP => CLK_I, Q => 
                           n_2684, QN => n2914);
   KEY_EXPAN0_reg_49_25_inst : FD1 port map( D => n6254, CP => CLK_I, Q => 
                           n_2685, QN => n2917);
   KEY_EXPAN0_reg_48_25_inst : FD1 port map( D => n6253, CP => CLK_I, Q => 
                           n_2686, QN => n2916);
   KEY_EXPAN0_reg_47_25_inst : FD1 port map( D => n6252, CP => CLK_I, Q => 
                           n_2687, QN => n2903);
   KEY_EXPAN0_reg_46_25_inst : FD1 port map( D => n6251, CP => CLK_I, Q => 
                           n_2688, QN => n2902);
   KEY_EXPAN0_reg_45_25_inst : FD1 port map( D => n6250, CP => CLK_I, Q => 
                           n_2689, QN => n2905);
   KEY_EXPAN0_reg_44_25_inst : FD1 port map( D => n6249, CP => CLK_I, Q => 
                           n_2690, QN => n2904);
   KEY_EXPAN0_reg_43_25_inst : FD1 port map( D => n6248, CP => CLK_I, Q => 
                           n_2691, QN => n2907);
   KEY_EXPAN0_reg_42_25_inst : FD1 port map( D => n6247, CP => CLK_I, Q => 
                           n_2692, QN => n2906);
   KEY_EXPAN0_reg_41_25_inst : FD1 port map( D => n6246, CP => CLK_I, Q => 
                           n_2693, QN => n2909);
   KEY_EXPAN0_reg_40_25_inst : FD1 port map( D => n6245, CP => CLK_I, Q => 
                           n_2694, QN => n2908);
   KEY_EXPAN0_reg_39_25_inst : FD1 port map( D => n6244, CP => CLK_I, Q => 
                           n_2695, QN => n2895);
   KEY_EXPAN0_reg_38_25_inst : FD1 port map( D => n6243, CP => CLK_I, Q => 
                           n_2696, QN => n2894);
   KEY_EXPAN0_reg_37_25_inst : FD1 port map( D => n6242, CP => CLK_I, Q => 
                           n_2697, QN => n2897);
   KEY_EXPAN0_reg_36_25_inst : FD1 port map( D => n6241, CP => CLK_I, Q => 
                           n_2698, QN => n2896);
   KEY_EXPAN0_reg_35_25_inst : FD1 port map( D => n6240, CP => CLK_I, Q => 
                           n_2699, QN => n2899);
   KEY_EXPAN0_reg_34_25_inst : FD1 port map( D => n6239, CP => CLK_I, Q => 
                           n_2700, QN => n2898);
   KEY_EXPAN0_reg_33_25_inst : FD1 port map( D => n6238, CP => CLK_I, Q => 
                           n_2701, QN => n2901);
   KEY_EXPAN0_reg_32_25_inst : FD1 port map( D => n6237, CP => CLK_I, Q => 
                           n_2702, QN => n2900);
   KEY_EXPAN0_reg_31_25_inst : FD1 port map( D => n6236, CP => CLK_I, Q => 
                           n_2703, QN => n2951);
   KEY_EXPAN0_reg_30_25_inst : FD1 port map( D => n6235, CP => CLK_I, Q => 
                           n_2704, QN => n2950);
   KEY_EXPAN0_reg_29_25_inst : FD1 port map( D => n6234, CP => CLK_I, Q => 
                           n_2705, QN => n2953);
   KEY_EXPAN0_reg_28_25_inst : FD1 port map( D => n6233, CP => CLK_I, Q => 
                           n_2706, QN => n2952);
   KEY_EXPAN0_reg_27_25_inst : FD1 port map( D => n6232, CP => CLK_I, Q => 
                           n_2707, QN => n2955);
   KEY_EXPAN0_reg_26_25_inst : FD1 port map( D => n6231, CP => CLK_I, Q => 
                           n_2708, QN => n2954);
   KEY_EXPAN0_reg_25_25_inst : FD1 port map( D => n6230, CP => CLK_I, Q => 
                           n_2709, QN => n2957);
   KEY_EXPAN0_reg_24_25_inst : FD1 port map( D => n6229, CP => CLK_I, Q => 
                           n_2710, QN => n2956);
   KEY_EXPAN0_reg_23_25_inst : FD1 port map( D => n6228, CP => CLK_I, Q => 
                           n_2711, QN => n2943);
   KEY_EXPAN0_reg_22_25_inst : FD1 port map( D => n6227, CP => CLK_I, Q => 
                           n_2712, QN => n2942);
   KEY_EXPAN0_reg_21_25_inst : FD1 port map( D => n6226, CP => CLK_I, Q => 
                           n_2713, QN => n2945);
   KEY_EXPAN0_reg_20_25_inst : FD1 port map( D => n6225, CP => CLK_I, Q => 
                           n_2714, QN => n2944);
   KEY_EXPAN0_reg_19_25_inst : FD1 port map( D => n6224, CP => CLK_I, Q => 
                           n_2715, QN => n2947);
   KEY_EXPAN0_reg_18_25_inst : FD1 port map( D => n6223, CP => CLK_I, Q => 
                           n_2716, QN => n2946);
   KEY_EXPAN0_reg_17_25_inst : FD1 port map( D => n6222, CP => CLK_I, Q => 
                           n_2717, QN => n2949);
   KEY_EXPAN0_reg_16_25_inst : FD1 port map( D => n6221, CP => CLK_I, Q => 
                           n_2718, QN => n2948);
   KEY_EXPAN0_reg_15_25_inst : FD1 port map( D => n6220, CP => CLK_I, Q => 
                           n_2719, QN => n2935);
   KEY_EXPAN0_reg_14_25_inst : FD1 port map( D => n6219, CP => CLK_I, Q => 
                           n_2720, QN => n2934);
   KEY_EXPAN0_reg_13_25_inst : FD1 port map( D => n6218, CP => CLK_I, Q => 
                           n_2721, QN => n2937);
   KEY_EXPAN0_reg_12_25_inst : FD1 port map( D => n6217, CP => CLK_I, Q => 
                           n_2722, QN => n2936);
   KEY_EXPAN0_reg_11_25_inst : FD1 port map( D => n6216, CP => CLK_I, Q => 
                           n_2723, QN => n2939);
   KEY_EXPAN0_reg_10_25_inst : FD1 port map( D => n6215, CP => CLK_I, Q => 
                           n_2724, QN => n2938);
   KEY_EXPAN0_reg_9_25_inst : FD1 port map( D => n6214, CP => CLK_I, Q => 
                           n_2725, QN => n2941);
   KEY_EXPAN0_reg_8_25_inst : FD1 port map( D => n6213, CP => CLK_I, Q => 
                           n_2726, QN => n2940);
   KEY_EXPAN0_reg_7_25_inst : FD1 port map( D => n6212, CP => CLK_I, Q => 
                           n_2727, QN => n2927);
   KEY_EXPAN0_reg_6_25_inst : FD1 port map( D => n6211, CP => CLK_I, Q => 
                           n_2728, QN => n2926);
   KEY_EXPAN0_reg_5_25_inst : FD1 port map( D => n6210, CP => CLK_I, Q => 
                           n_2729, QN => n2929);
   KEY_EXPAN0_reg_4_25_inst : FD1 port map( D => n6209, CP => CLK_I, Q => 
                           n_2730, QN => n2928);
   KEY_EXPAN0_reg_3_25_inst : FD1 port map( D => n6208, CP => CLK_I, Q => 
                           n_2731, QN => n2931);
   KEY_EXPAN0_reg_2_25_inst : FD1 port map( D => n6207, CP => CLK_I, Q => 
                           n_2732, QN => n2930);
   KEY_EXPAN0_reg_1_25_inst : FD1 port map( D => n6206, CP => CLK_I, Q => 
                           n_2733, QN => n2933);
   KEY_EXPAN0_reg_0_25_inst : FD1 port map( D => n6205, CP => CLK_I, Q => 
                           n_2734, QN => n2932);
   v_KEY_COL_OUT0_reg_25_inst : FD1 port map( D => n4570, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_25_port, QN => n1989);
   v_TEMP_VECTOR_reg_17_inst : FD1 port map( D => n6692, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_17_port, QN => n_2735);
   KEY_EXPAN0_reg_63_17_inst : FD1 port map( D => n5756, CP => CLK_I, Q => 
                           n_2736, QN => n2855);
   KEY_EXPAN0_reg_62_17_inst : FD1 port map( D => n5755, CP => CLK_I, Q => 
                           n_2737, QN => n2854);
   KEY_EXPAN0_reg_61_17_inst : FD1 port map( D => n5754, CP => CLK_I, Q => 
                           n_2738, QN => n2857);
   KEY_EXPAN0_reg_60_17_inst : FD1 port map( D => n5753, CP => CLK_I, Q => 
                           n_2739, QN => n2856);
   KEY_EXPAN0_reg_59_17_inst : FD1 port map( D => n5752, CP => CLK_I, Q => 
                           n_2740, QN => n2859);
   KEY_EXPAN0_reg_58_17_inst : FD1 port map( D => n5751, CP => CLK_I, Q => 
                           n_2741, QN => n2858);
   KEY_EXPAN0_reg_57_17_inst : FD1 port map( D => n5750, CP => CLK_I, Q => 
                           n_2742, QN => n2861);
   KEY_EXPAN0_reg_56_17_inst : FD1 port map( D => n5749, CP => CLK_I, Q => 
                           n_2743, QN => n2860);
   KEY_EXPAN0_reg_55_17_inst : FD1 port map( D => n5748, CP => CLK_I, Q => 
                           n_2744, QN => n2847);
   KEY_EXPAN0_reg_54_17_inst : FD1 port map( D => n5747, CP => CLK_I, Q => 
                           n_2745, QN => n2846);
   KEY_EXPAN0_reg_53_17_inst : FD1 port map( D => n5746, CP => CLK_I, Q => 
                           n_2746, QN => n2849);
   KEY_EXPAN0_reg_52_17_inst : FD1 port map( D => n5745, CP => CLK_I, Q => 
                           n_2747, QN => n2848);
   KEY_EXPAN0_reg_51_17_inst : FD1 port map( D => n5744, CP => CLK_I, Q => 
                           n_2748, QN => n2851);
   KEY_EXPAN0_reg_50_17_inst : FD1 port map( D => n5743, CP => CLK_I, Q => 
                           n_2749, QN => n2850);
   KEY_EXPAN0_reg_49_17_inst : FD1 port map( D => n5742, CP => CLK_I, Q => 
                           n_2750, QN => n2853);
   KEY_EXPAN0_reg_48_17_inst : FD1 port map( D => n5741, CP => CLK_I, Q => 
                           n_2751, QN => n2852);
   KEY_EXPAN0_reg_47_17_inst : FD1 port map( D => n5740, CP => CLK_I, Q => 
                           n_2752, QN => n2839);
   KEY_EXPAN0_reg_46_17_inst : FD1 port map( D => n5739, CP => CLK_I, Q => 
                           n_2753, QN => n2838);
   KEY_EXPAN0_reg_45_17_inst : FD1 port map( D => n5738, CP => CLK_I, Q => 
                           n_2754, QN => n2841);
   KEY_EXPAN0_reg_44_17_inst : FD1 port map( D => n5737, CP => CLK_I, Q => 
                           n_2755, QN => n2840);
   KEY_EXPAN0_reg_43_17_inst : FD1 port map( D => n5736, CP => CLK_I, Q => 
                           n_2756, QN => n2843);
   KEY_EXPAN0_reg_42_17_inst : FD1 port map( D => n5735, CP => CLK_I, Q => 
                           n_2757, QN => n2842);
   KEY_EXPAN0_reg_41_17_inst : FD1 port map( D => n5734, CP => CLK_I, Q => 
                           n_2758, QN => n2845);
   KEY_EXPAN0_reg_40_17_inst : FD1 port map( D => n5733, CP => CLK_I, Q => 
                           n_2759, QN => n2844);
   KEY_EXPAN0_reg_39_17_inst : FD1 port map( D => n5732, CP => CLK_I, Q => 
                           n_2760, QN => n2831);
   KEY_EXPAN0_reg_38_17_inst : FD1 port map( D => n5731, CP => CLK_I, Q => 
                           n_2761, QN => n2830);
   KEY_EXPAN0_reg_37_17_inst : FD1 port map( D => n5730, CP => CLK_I, Q => 
                           n_2762, QN => n2833);
   KEY_EXPAN0_reg_36_17_inst : FD1 port map( D => n5729, CP => CLK_I, Q => 
                           n_2763, QN => n2832);
   KEY_EXPAN0_reg_35_17_inst : FD1 port map( D => n5728, CP => CLK_I, Q => 
                           n_2764, QN => n2835);
   KEY_EXPAN0_reg_34_17_inst : FD1 port map( D => n5727, CP => CLK_I, Q => 
                           n_2765, QN => n2834);
   KEY_EXPAN0_reg_33_17_inst : FD1 port map( D => n5726, CP => CLK_I, Q => 
                           n_2766, QN => n2837);
   KEY_EXPAN0_reg_32_17_inst : FD1 port map( D => n5725, CP => CLK_I, Q => 
                           n_2767, QN => n2836);
   KEY_EXPAN0_reg_31_17_inst : FD1 port map( D => n5724, CP => CLK_I, Q => 
                           n_2768, QN => n2887);
   KEY_EXPAN0_reg_30_17_inst : FD1 port map( D => n5723, CP => CLK_I, Q => 
                           n_2769, QN => n2886);
   KEY_EXPAN0_reg_29_17_inst : FD1 port map( D => n5722, CP => CLK_I, Q => 
                           n_2770, QN => n2889);
   KEY_EXPAN0_reg_28_17_inst : FD1 port map( D => n5721, CP => CLK_I, Q => 
                           n_2771, QN => n2888);
   KEY_EXPAN0_reg_27_17_inst : FD1 port map( D => n5720, CP => CLK_I, Q => 
                           n_2772, QN => n2891);
   KEY_EXPAN0_reg_26_17_inst : FD1 port map( D => n5719, CP => CLK_I, Q => 
                           n_2773, QN => n2890);
   KEY_EXPAN0_reg_25_17_inst : FD1 port map( D => n5718, CP => CLK_I, Q => 
                           n_2774, QN => n2893);
   KEY_EXPAN0_reg_24_17_inst : FD1 port map( D => n5717, CP => CLK_I, Q => 
                           n_2775, QN => n2892);
   KEY_EXPAN0_reg_23_17_inst : FD1 port map( D => n5716, CP => CLK_I, Q => 
                           n_2776, QN => n2879);
   KEY_EXPAN0_reg_22_17_inst : FD1 port map( D => n5715, CP => CLK_I, Q => 
                           n_2777, QN => n2878);
   KEY_EXPAN0_reg_21_17_inst : FD1 port map( D => n5714, CP => CLK_I, Q => 
                           n_2778, QN => n2881);
   KEY_EXPAN0_reg_20_17_inst : FD1 port map( D => n5713, CP => CLK_I, Q => 
                           n_2779, QN => n2880);
   KEY_EXPAN0_reg_19_17_inst : FD1 port map( D => n5712, CP => CLK_I, Q => 
                           n_2780, QN => n2883);
   KEY_EXPAN0_reg_18_17_inst : FD1 port map( D => n5711, CP => CLK_I, Q => 
                           n_2781, QN => n2882);
   KEY_EXPAN0_reg_17_17_inst : FD1 port map( D => n5710, CP => CLK_I, Q => 
                           n_2782, QN => n2885);
   KEY_EXPAN0_reg_16_17_inst : FD1 port map( D => n5709, CP => CLK_I, Q => 
                           n_2783, QN => n2884);
   KEY_EXPAN0_reg_15_17_inst : FD1 port map( D => n5708, CP => CLK_I, Q => 
                           n_2784, QN => n2871);
   KEY_EXPAN0_reg_14_17_inst : FD1 port map( D => n5707, CP => CLK_I, Q => 
                           n_2785, QN => n2870);
   KEY_EXPAN0_reg_13_17_inst : FD1 port map( D => n5706, CP => CLK_I, Q => 
                           n_2786, QN => n2873);
   KEY_EXPAN0_reg_12_17_inst : FD1 port map( D => n5705, CP => CLK_I, Q => 
                           n_2787, QN => n2872);
   KEY_EXPAN0_reg_11_17_inst : FD1 port map( D => n5704, CP => CLK_I, Q => 
                           n_2788, QN => n2875);
   KEY_EXPAN0_reg_10_17_inst : FD1 port map( D => n5703, CP => CLK_I, Q => 
                           n_2789, QN => n2874);
   KEY_EXPAN0_reg_9_17_inst : FD1 port map( D => n5702, CP => CLK_I, Q => 
                           n_2790, QN => n2877);
   KEY_EXPAN0_reg_8_17_inst : FD1 port map( D => n5701, CP => CLK_I, Q => 
                           n_2791, QN => n2876);
   KEY_EXPAN0_reg_7_17_inst : FD1 port map( D => n5700, CP => CLK_I, Q => 
                           n_2792, QN => n2863);
   KEY_EXPAN0_reg_6_17_inst : FD1 port map( D => n5699, CP => CLK_I, Q => 
                           n_2793, QN => n2862);
   KEY_EXPAN0_reg_5_17_inst : FD1 port map( D => n5698, CP => CLK_I, Q => 
                           n_2794, QN => n2865);
   KEY_EXPAN0_reg_4_17_inst : FD1 port map( D => n5697, CP => CLK_I, Q => 
                           n_2795, QN => n2864);
   KEY_EXPAN0_reg_3_17_inst : FD1 port map( D => n5696, CP => CLK_I, Q => 
                           n_2796, QN => n2867);
   KEY_EXPAN0_reg_2_17_inst : FD1 port map( D => n5695, CP => CLK_I, Q => 
                           n_2797, QN => n2866);
   KEY_EXPAN0_reg_1_17_inst : FD1 port map( D => n5694, CP => CLK_I, Q => 
                           n_2798, QN => n2869);
   KEY_EXPAN0_reg_0_17_inst : FD1 port map( D => n5693, CP => CLK_I, Q => 
                           n_2799, QN => n2868);
   v_KEY_COL_OUT0_reg_17_inst : FD1 port map( D => n4569, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_17_port, QN => n1949);
   v_TEMP_VECTOR_reg_9_inst : FD1 port map( D => n6700, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_9_port, QN => n_2800);
   KEY_EXPAN0_reg_63_9_inst : FD1 port map( D => n5244, CP => CLK_I, Q => 
                           n_2801, QN => n2791);
   KEY_EXPAN0_reg_62_9_inst : FD1 port map( D => n5243, CP => CLK_I, Q => 
                           n_2802, QN => n2790);
   KEY_EXPAN0_reg_61_9_inst : FD1 port map( D => n5242, CP => CLK_I, Q => 
                           n_2803, QN => n2793);
   KEY_EXPAN0_reg_60_9_inst : FD1 port map( D => n5241, CP => CLK_I, Q => 
                           n_2804, QN => n2792);
   KEY_EXPAN0_reg_59_9_inst : FD1 port map( D => n5240, CP => CLK_I, Q => 
                           n_2805, QN => n2795);
   KEY_EXPAN0_reg_58_9_inst : FD1 port map( D => n5239, CP => CLK_I, Q => 
                           n_2806, QN => n2794);
   KEY_EXPAN0_reg_57_9_inst : FD1 port map( D => n5238, CP => CLK_I, Q => 
                           n_2807, QN => n2797);
   KEY_EXPAN0_reg_56_9_inst : FD1 port map( D => n5237, CP => CLK_I, Q => 
                           n_2808, QN => n2796);
   KEY_EXPAN0_reg_55_9_inst : FD1 port map( D => n5236, CP => CLK_I, Q => 
                           n_2809, QN => n2783);
   KEY_EXPAN0_reg_54_9_inst : FD1 port map( D => n5235, CP => CLK_I, Q => 
                           n_2810, QN => n2782);
   KEY_EXPAN0_reg_53_9_inst : FD1 port map( D => n5234, CP => CLK_I, Q => 
                           n_2811, QN => n2785);
   KEY_EXPAN0_reg_52_9_inst : FD1 port map( D => n5233, CP => CLK_I, Q => 
                           n_2812, QN => n2784);
   KEY_EXPAN0_reg_51_9_inst : FD1 port map( D => n5232, CP => CLK_I, Q => 
                           n_2813, QN => n2787);
   KEY_EXPAN0_reg_50_9_inst : FD1 port map( D => n5231, CP => CLK_I, Q => 
                           n_2814, QN => n2786);
   KEY_EXPAN0_reg_49_9_inst : FD1 port map( D => n5230, CP => CLK_I, Q => 
                           n_2815, QN => n2789);
   KEY_EXPAN0_reg_48_9_inst : FD1 port map( D => n5229, CP => CLK_I, Q => 
                           n_2816, QN => n2788);
   KEY_EXPAN0_reg_47_9_inst : FD1 port map( D => n5228, CP => CLK_I, Q => 
                           n_2817, QN => n2775);
   KEY_EXPAN0_reg_46_9_inst : FD1 port map( D => n5227, CP => CLK_I, Q => 
                           n_2818, QN => n2774);
   KEY_EXPAN0_reg_45_9_inst : FD1 port map( D => n5226, CP => CLK_I, Q => 
                           n_2819, QN => n2777);
   KEY_EXPAN0_reg_44_9_inst : FD1 port map( D => n5225, CP => CLK_I, Q => 
                           n_2820, QN => n2776);
   KEY_EXPAN0_reg_43_9_inst : FD1 port map( D => n5224, CP => CLK_I, Q => 
                           n_2821, QN => n2779);
   KEY_EXPAN0_reg_42_9_inst : FD1 port map( D => n5223, CP => CLK_I, Q => 
                           n_2822, QN => n2778);
   KEY_EXPAN0_reg_41_9_inst : FD1 port map( D => n5222, CP => CLK_I, Q => 
                           n_2823, QN => n2781);
   KEY_EXPAN0_reg_40_9_inst : FD1 port map( D => n5221, CP => CLK_I, Q => 
                           n_2824, QN => n2780);
   KEY_EXPAN0_reg_39_9_inst : FD1 port map( D => n5220, CP => CLK_I, Q => 
                           n_2825, QN => n2767);
   KEY_EXPAN0_reg_38_9_inst : FD1 port map( D => n5219, CP => CLK_I, Q => 
                           n_2826, QN => n2766);
   KEY_EXPAN0_reg_37_9_inst : FD1 port map( D => n5218, CP => CLK_I, Q => 
                           n_2827, QN => n2769);
   KEY_EXPAN0_reg_36_9_inst : FD1 port map( D => n5217, CP => CLK_I, Q => 
                           n_2828, QN => n2768);
   KEY_EXPAN0_reg_35_9_inst : FD1 port map( D => n5216, CP => CLK_I, Q => 
                           n_2829, QN => n2771);
   KEY_EXPAN0_reg_34_9_inst : FD1 port map( D => n5215, CP => CLK_I, Q => 
                           n_2830, QN => n2770);
   KEY_EXPAN0_reg_33_9_inst : FD1 port map( D => n5214, CP => CLK_I, Q => 
                           n_2831, QN => n2773);
   KEY_EXPAN0_reg_32_9_inst : FD1 port map( D => n5213, CP => CLK_I, Q => 
                           n_2832, QN => n2772);
   KEY_EXPAN0_reg_31_9_inst : FD1 port map( D => n5212, CP => CLK_I, Q => 
                           n_2833, QN => n2823);
   KEY_EXPAN0_reg_30_9_inst : FD1 port map( D => n5211, CP => CLK_I, Q => 
                           n_2834, QN => n2822);
   KEY_EXPAN0_reg_29_9_inst : FD1 port map( D => n5210, CP => CLK_I, Q => 
                           n_2835, QN => n2825);
   KEY_EXPAN0_reg_28_9_inst : FD1 port map( D => n5209, CP => CLK_I, Q => 
                           n_2836, QN => n2824);
   KEY_EXPAN0_reg_27_9_inst : FD1 port map( D => n5208, CP => CLK_I, Q => 
                           n_2837, QN => n2827);
   KEY_EXPAN0_reg_26_9_inst : FD1 port map( D => n5207, CP => CLK_I, Q => 
                           n_2838, QN => n2826);
   KEY_EXPAN0_reg_25_9_inst : FD1 port map( D => n5206, CP => CLK_I, Q => 
                           n_2839, QN => n2829);
   KEY_EXPAN0_reg_24_9_inst : FD1 port map( D => n5205, CP => CLK_I, Q => 
                           n_2840, QN => n2828);
   KEY_EXPAN0_reg_23_9_inst : FD1 port map( D => n5204, CP => CLK_I, Q => 
                           n_2841, QN => n2815);
   KEY_EXPAN0_reg_22_9_inst : FD1 port map( D => n5203, CP => CLK_I, Q => 
                           n_2842, QN => n2814);
   KEY_EXPAN0_reg_21_9_inst : FD1 port map( D => n5202, CP => CLK_I, Q => 
                           n_2843, QN => n2817);
   KEY_EXPAN0_reg_20_9_inst : FD1 port map( D => n5201, CP => CLK_I, Q => 
                           n_2844, QN => n2816);
   KEY_EXPAN0_reg_19_9_inst : FD1 port map( D => n5200, CP => CLK_I, Q => 
                           n_2845, QN => n2819);
   KEY_EXPAN0_reg_18_9_inst : FD1 port map( D => n5199, CP => CLK_I, Q => 
                           n_2846, QN => n2818);
   KEY_EXPAN0_reg_17_9_inst : FD1 port map( D => n5198, CP => CLK_I, Q => 
                           n_2847, QN => n2821);
   KEY_EXPAN0_reg_16_9_inst : FD1 port map( D => n5197, CP => CLK_I, Q => 
                           n_2848, QN => n2820);
   KEY_EXPAN0_reg_15_9_inst : FD1 port map( D => n5196, CP => CLK_I, Q => 
                           n_2849, QN => n2807);
   KEY_EXPAN0_reg_14_9_inst : FD1 port map( D => n5195, CP => CLK_I, Q => 
                           n_2850, QN => n2806);
   KEY_EXPAN0_reg_13_9_inst : FD1 port map( D => n5194, CP => CLK_I, Q => 
                           n_2851, QN => n2809);
   KEY_EXPAN0_reg_12_9_inst : FD1 port map( D => n5193, CP => CLK_I, Q => 
                           n_2852, QN => n2808);
   KEY_EXPAN0_reg_11_9_inst : FD1 port map( D => n5192, CP => CLK_I, Q => 
                           n_2853, QN => n2811);
   KEY_EXPAN0_reg_10_9_inst : FD1 port map( D => n5191, CP => CLK_I, Q => 
                           n_2854, QN => n2810);
   KEY_EXPAN0_reg_9_9_inst : FD1 port map( D => n5190, CP => CLK_I, Q => n_2855
                           , QN => n2813);
   KEY_EXPAN0_reg_8_9_inst : FD1 port map( D => n5189, CP => CLK_I, Q => n_2856
                           , QN => n2812);
   KEY_EXPAN0_reg_7_9_inst : FD1 port map( D => n5188, CP => CLK_I, Q => n_2857
                           , QN => n2799);
   KEY_EXPAN0_reg_6_9_inst : FD1 port map( D => n5187, CP => CLK_I, Q => n_2858
                           , QN => n2798);
   KEY_EXPAN0_reg_5_9_inst : FD1 port map( D => n5186, CP => CLK_I, Q => n_2859
                           , QN => n2801);
   KEY_EXPAN0_reg_4_9_inst : FD1 port map( D => n5185, CP => CLK_I, Q => n_2860
                           , QN => n2800);
   KEY_EXPAN0_reg_3_9_inst : FD1 port map( D => n5184, CP => CLK_I, Q => n_2861
                           , QN => n2803);
   KEY_EXPAN0_reg_2_9_inst : FD1 port map( D => n5183, CP => CLK_I, Q => n_2862
                           , QN => n2802);
   KEY_EXPAN0_reg_1_9_inst : FD1 port map( D => n5182, CP => CLK_I, Q => n_2863
                           , QN => n2805);
   KEY_EXPAN0_reg_0_9_inst : FD1 port map( D => n5181, CP => CLK_I, Q => n_2864
                           , QN => n2804);
   v_KEY_COL_OUT0_reg_9_inst : FD1 port map( D => n4568, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_9_port, QN => n1974);
   v_TEMP_VECTOR_reg_0_inst : FD1 port map( D => n6709, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_0_port, QN => n2103);
   KEY_EXPAN0_reg_63_0_inst : FD1 port map( D => n4668, CP => CLK_I, Q => 
                           n_2865, QN => n2727);
   KEY_EXPAN0_reg_62_0_inst : FD1 port map( D => n4667, CP => CLK_I, Q => 
                           n_2866, QN => n2726);
   KEY_EXPAN0_reg_61_0_inst : FD1 port map( D => n4666, CP => CLK_I, Q => 
                           n_2867, QN => n2729);
   KEY_EXPAN0_reg_60_0_inst : FD1 port map( D => n4665, CP => CLK_I, Q => 
                           n_2868, QN => n2728);
   KEY_EXPAN0_reg_59_0_inst : FD1 port map( D => n4664, CP => CLK_I, Q => 
                           n_2869, QN => n2731);
   KEY_EXPAN0_reg_58_0_inst : FD1 port map( D => n4663, CP => CLK_I, Q => 
                           n_2870, QN => n2730);
   KEY_EXPAN0_reg_57_0_inst : FD1 port map( D => n4662, CP => CLK_I, Q => 
                           n_2871, QN => n2733);
   KEY_EXPAN0_reg_56_0_inst : FD1 port map( D => n4661, CP => CLK_I, Q => 
                           n_2872, QN => n2732);
   KEY_EXPAN0_reg_55_0_inst : FD1 port map( D => n4660, CP => CLK_I, Q => 
                           n_2873, QN => n2719);
   KEY_EXPAN0_reg_54_0_inst : FD1 port map( D => n4659, CP => CLK_I, Q => 
                           n_2874, QN => n2718);
   KEY_EXPAN0_reg_53_0_inst : FD1 port map( D => n4658, CP => CLK_I, Q => 
                           n_2875, QN => n2721);
   KEY_EXPAN0_reg_52_0_inst : FD1 port map( D => n4657, CP => CLK_I, Q => 
                           n_2876, QN => n2720);
   KEY_EXPAN0_reg_51_0_inst : FD1 port map( D => n4656, CP => CLK_I, Q => 
                           n_2877, QN => n2723);
   KEY_EXPAN0_reg_50_0_inst : FD1 port map( D => n4655, CP => CLK_I, Q => 
                           n_2878, QN => n2722);
   KEY_EXPAN0_reg_49_0_inst : FD1 port map( D => n4654, CP => CLK_I, Q => 
                           n_2879, QN => n2725);
   KEY_EXPAN0_reg_48_0_inst : FD1 port map( D => n4653, CP => CLK_I, Q => 
                           n_2880, QN => n2724);
   KEY_EXPAN0_reg_47_0_inst : FD1 port map( D => n4652, CP => CLK_I, Q => 
                           n_2881, QN => n2711);
   KEY_EXPAN0_reg_46_0_inst : FD1 port map( D => n4651, CP => CLK_I, Q => 
                           n_2882, QN => n2710);
   KEY_EXPAN0_reg_45_0_inst : FD1 port map( D => n4650, CP => CLK_I, Q => 
                           n_2883, QN => n2713);
   KEY_EXPAN0_reg_44_0_inst : FD1 port map( D => n4649, CP => CLK_I, Q => 
                           n_2884, QN => n2712);
   KEY_EXPAN0_reg_43_0_inst : FD1 port map( D => n4648, CP => CLK_I, Q => 
                           n_2885, QN => n2715);
   KEY_EXPAN0_reg_42_0_inst : FD1 port map( D => n4647, CP => CLK_I, Q => 
                           n_2886, QN => n2714);
   KEY_EXPAN0_reg_41_0_inst : FD1 port map( D => n4646, CP => CLK_I, Q => 
                           n_2887, QN => n2717);
   KEY_EXPAN0_reg_40_0_inst : FD1 port map( D => n4645, CP => CLK_I, Q => 
                           n_2888, QN => n2716);
   KEY_EXPAN0_reg_39_0_inst : FD1 port map( D => n4644, CP => CLK_I, Q => 
                           n_2889, QN => n2703);
   KEY_EXPAN0_reg_38_0_inst : FD1 port map( D => n4643, CP => CLK_I, Q => 
                           n_2890, QN => n2702);
   KEY_EXPAN0_reg_37_0_inst : FD1 port map( D => n4642, CP => CLK_I, Q => 
                           n_2891, QN => n2705);
   KEY_EXPAN0_reg_36_0_inst : FD1 port map( D => n4641, CP => CLK_I, Q => 
                           n_2892, QN => n2704);
   KEY_EXPAN0_reg_35_0_inst : FD1 port map( D => n4640, CP => CLK_I, Q => 
                           n_2893, QN => n2707);
   KEY_EXPAN0_reg_34_0_inst : FD1 port map( D => n4639, CP => CLK_I, Q => 
                           n_2894, QN => n2706);
   KEY_EXPAN0_reg_33_0_inst : FD1 port map( D => n4638, CP => CLK_I, Q => 
                           n_2895, QN => n2709);
   KEY_EXPAN0_reg_32_0_inst : FD1 port map( D => n4637, CP => CLK_I, Q => 
                           n_2896, QN => n2708);
   KEY_EXPAN0_reg_31_0_inst : FD1 port map( D => n4636, CP => CLK_I, Q => 
                           n_2897, QN => n2759);
   KEY_EXPAN0_reg_30_0_inst : FD1 port map( D => n4635, CP => CLK_I, Q => 
                           n_2898, QN => n2758);
   KEY_EXPAN0_reg_29_0_inst : FD1 port map( D => n4634, CP => CLK_I, Q => 
                           n_2899, QN => n2761);
   KEY_EXPAN0_reg_28_0_inst : FD1 port map( D => n4633, CP => CLK_I, Q => 
                           n_2900, QN => n2760);
   KEY_EXPAN0_reg_27_0_inst : FD1 port map( D => n4632, CP => CLK_I, Q => 
                           n_2901, QN => n2763);
   KEY_EXPAN0_reg_26_0_inst : FD1 port map( D => n4631, CP => CLK_I, Q => 
                           n_2902, QN => n2762);
   KEY_EXPAN0_reg_25_0_inst : FD1 port map( D => n4630, CP => CLK_I, Q => 
                           n_2903, QN => n2765);
   KEY_EXPAN0_reg_24_0_inst : FD1 port map( D => n4629, CP => CLK_I, Q => 
                           n_2904, QN => n2764);
   KEY_EXPAN0_reg_23_0_inst : FD1 port map( D => n4628, CP => CLK_I, Q => 
                           n_2905, QN => n2751);
   KEY_EXPAN0_reg_22_0_inst : FD1 port map( D => n4627, CP => CLK_I, Q => 
                           n_2906, QN => n2750);
   KEY_EXPAN0_reg_21_0_inst : FD1 port map( D => n4626, CP => CLK_I, Q => 
                           n_2907, QN => n2753);
   KEY_EXPAN0_reg_20_0_inst : FD1 port map( D => n4625, CP => CLK_I, Q => 
                           n_2908, QN => n2752);
   KEY_EXPAN0_reg_19_0_inst : FD1 port map( D => n4624, CP => CLK_I, Q => 
                           n_2909, QN => n2755);
   KEY_EXPAN0_reg_18_0_inst : FD1 port map( D => n4623, CP => CLK_I, Q => 
                           n_2910, QN => n2754);
   KEY_EXPAN0_reg_17_0_inst : FD1 port map( D => n4622, CP => CLK_I, Q => 
                           n_2911, QN => n2757);
   KEY_EXPAN0_reg_16_0_inst : FD1 port map( D => n4621, CP => CLK_I, Q => 
                           n_2912, QN => n2756);
   KEY_EXPAN0_reg_15_0_inst : FD1 port map( D => n4620, CP => CLK_I, Q => 
                           n_2913, QN => n2743);
   KEY_EXPAN0_reg_14_0_inst : FD1 port map( D => n4619, CP => CLK_I, Q => 
                           n_2914, QN => n2742);
   KEY_EXPAN0_reg_13_0_inst : FD1 port map( D => n4618, CP => CLK_I, Q => 
                           n_2915, QN => n2745);
   KEY_EXPAN0_reg_12_0_inst : FD1 port map( D => n4617, CP => CLK_I, Q => 
                           n_2916, QN => n2744);
   KEY_EXPAN0_reg_11_0_inst : FD1 port map( D => n4616, CP => CLK_I, Q => 
                           n_2917, QN => n2747);
   KEY_EXPAN0_reg_10_0_inst : FD1 port map( D => n4615, CP => CLK_I, Q => 
                           n_2918, QN => n2746);
   KEY_EXPAN0_reg_9_0_inst : FD1 port map( D => n4614, CP => CLK_I, Q => n_2919
                           , QN => n2749);
   KEY_EXPAN0_reg_8_0_inst : FD1 port map( D => n4613, CP => CLK_I, Q => n_2920
                           , QN => n2748);
   KEY_EXPAN0_reg_7_0_inst : FD1 port map( D => n4612, CP => CLK_I, Q => n_2921
                           , QN => n2735);
   KEY_EXPAN0_reg_6_0_inst : FD1 port map( D => n4611, CP => CLK_I, Q => n_2922
                           , QN => n2734);
   KEY_EXPAN0_reg_5_0_inst : FD1 port map( D => n4610, CP => CLK_I, Q => n_2923
                           , QN => n2737);
   KEY_EXPAN0_reg_4_0_inst : FD1 port map( D => n4609, CP => CLK_I, Q => n_2924
                           , QN => n2736);
   KEY_EXPAN0_reg_3_0_inst : FD1 port map( D => n4608, CP => CLK_I, Q => n_2925
                           , QN => n2739);
   KEY_EXPAN0_reg_2_0_inst : FD1 port map( D => n4607, CP => CLK_I, Q => n_2926
                           , QN => n2738);
   KEY_EXPAN0_reg_1_0_inst : FD1 port map( D => n4606, CP => CLK_I, Q => n_2927
                           , QN => n2741);
   KEY_EXPAN0_reg_0_0_inst : FD1 port map( D => n4605, CP => CLK_I, Q => n_2928
                           , QN => n2740);
   v_KEY_COL_OUT0_reg_0_inst : FD1 port map( D => n4567, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_0_port, QN => n1981);
   v_TEMP_VECTOR_reg_24_inst : FD1 port map( D => n6685, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_24_port, QN => n_2929);
   KEY_EXPAN0_reg_63_24_inst : FD1 port map( D => n6204, CP => CLK_I, Q => 
                           n_2930, QN => n2663);
   KEY_EXPAN0_reg_62_24_inst : FD1 port map( D => n6203, CP => CLK_I, Q => 
                           n_2931, QN => n2662);
   KEY_EXPAN0_reg_61_24_inst : FD1 port map( D => n6202, CP => CLK_I, Q => 
                           n_2932, QN => n2665);
   KEY_EXPAN0_reg_60_24_inst : FD1 port map( D => n6201, CP => CLK_I, Q => 
                           n_2933, QN => n2664);
   KEY_EXPAN0_reg_59_24_inst : FD1 port map( D => n6200, CP => CLK_I, Q => 
                           n_2934, QN => n2667);
   KEY_EXPAN0_reg_58_24_inst : FD1 port map( D => n6199, CP => CLK_I, Q => 
                           n_2935, QN => n2666);
   KEY_EXPAN0_reg_57_24_inst : FD1 port map( D => n6198, CP => CLK_I, Q => 
                           n_2936, QN => n2669);
   KEY_EXPAN0_reg_56_24_inst : FD1 port map( D => n6197, CP => CLK_I, Q => 
                           n_2937, QN => n2668);
   KEY_EXPAN0_reg_55_24_inst : FD1 port map( D => n6196, CP => CLK_I, Q => 
                           n_2938, QN => n2655);
   KEY_EXPAN0_reg_54_24_inst : FD1 port map( D => n6195, CP => CLK_I, Q => 
                           n_2939, QN => n2654);
   KEY_EXPAN0_reg_53_24_inst : FD1 port map( D => n6194, CP => CLK_I, Q => 
                           n_2940, QN => n2657);
   KEY_EXPAN0_reg_52_24_inst : FD1 port map( D => n6193, CP => CLK_I, Q => 
                           n_2941, QN => n2656);
   KEY_EXPAN0_reg_51_24_inst : FD1 port map( D => n6192, CP => CLK_I, Q => 
                           n_2942, QN => n2659);
   KEY_EXPAN0_reg_50_24_inst : FD1 port map( D => n6191, CP => CLK_I, Q => 
                           n_2943, QN => n2658);
   KEY_EXPAN0_reg_49_24_inst : FD1 port map( D => n6190, CP => CLK_I, Q => 
                           n_2944, QN => n2661);
   KEY_EXPAN0_reg_48_24_inst : FD1 port map( D => n6189, CP => CLK_I, Q => 
                           n_2945, QN => n2660);
   KEY_EXPAN0_reg_47_24_inst : FD1 port map( D => n6188, CP => CLK_I, Q => 
                           n_2946, QN => n2647);
   KEY_EXPAN0_reg_46_24_inst : FD1 port map( D => n6187, CP => CLK_I, Q => 
                           n_2947, QN => n2646);
   KEY_EXPAN0_reg_45_24_inst : FD1 port map( D => n6186, CP => CLK_I, Q => 
                           n_2948, QN => n2649);
   KEY_EXPAN0_reg_44_24_inst : FD1 port map( D => n6185, CP => CLK_I, Q => 
                           n_2949, QN => n2648);
   KEY_EXPAN0_reg_43_24_inst : FD1 port map( D => n6184, CP => CLK_I, Q => 
                           n_2950, QN => n2651);
   KEY_EXPAN0_reg_42_24_inst : FD1 port map( D => n6183, CP => CLK_I, Q => 
                           n_2951, QN => n2650);
   KEY_EXPAN0_reg_41_24_inst : FD1 port map( D => n6182, CP => CLK_I, Q => 
                           n_2952, QN => n2653);
   KEY_EXPAN0_reg_40_24_inst : FD1 port map( D => n6181, CP => CLK_I, Q => 
                           n_2953, QN => n2652);
   KEY_EXPAN0_reg_39_24_inst : FD1 port map( D => n6180, CP => CLK_I, Q => 
                           n_2954, QN => n2639);
   KEY_EXPAN0_reg_38_24_inst : FD1 port map( D => n6179, CP => CLK_I, Q => 
                           n_2955, QN => n2638);
   KEY_EXPAN0_reg_37_24_inst : FD1 port map( D => n6178, CP => CLK_I, Q => 
                           n_2956, QN => n2641);
   KEY_EXPAN0_reg_36_24_inst : FD1 port map( D => n6177, CP => CLK_I, Q => 
                           n_2957, QN => n2640);
   KEY_EXPAN0_reg_35_24_inst : FD1 port map( D => n6176, CP => CLK_I, Q => 
                           n_2958, QN => n2643);
   KEY_EXPAN0_reg_34_24_inst : FD1 port map( D => n6175, CP => CLK_I, Q => 
                           n_2959, QN => n2642);
   KEY_EXPAN0_reg_33_24_inst : FD1 port map( D => n6174, CP => CLK_I, Q => 
                           n_2960, QN => n2645);
   KEY_EXPAN0_reg_32_24_inst : FD1 port map( D => n6173, CP => CLK_I, Q => 
                           n_2961, QN => n2644);
   KEY_EXPAN0_reg_31_24_inst : FD1 port map( D => n6172, CP => CLK_I, Q => 
                           n_2962, QN => n2695);
   KEY_EXPAN0_reg_30_24_inst : FD1 port map( D => n6171, CP => CLK_I, Q => 
                           n_2963, QN => n2694);
   KEY_EXPAN0_reg_29_24_inst : FD1 port map( D => n6170, CP => CLK_I, Q => 
                           n_2964, QN => n2697);
   KEY_EXPAN0_reg_28_24_inst : FD1 port map( D => n6169, CP => CLK_I, Q => 
                           n_2965, QN => n2696);
   KEY_EXPAN0_reg_27_24_inst : FD1 port map( D => n6168, CP => CLK_I, Q => 
                           n_2966, QN => n2699);
   KEY_EXPAN0_reg_26_24_inst : FD1 port map( D => n6167, CP => CLK_I, Q => 
                           n_2967, QN => n2698);
   KEY_EXPAN0_reg_25_24_inst : FD1 port map( D => n6166, CP => CLK_I, Q => 
                           n_2968, QN => n2701);
   KEY_EXPAN0_reg_24_24_inst : FD1 port map( D => n6165, CP => CLK_I, Q => 
                           n_2969, QN => n2700);
   KEY_EXPAN0_reg_23_24_inst : FD1 port map( D => n6164, CP => CLK_I, Q => 
                           n_2970, QN => n2687);
   KEY_EXPAN0_reg_22_24_inst : FD1 port map( D => n6163, CP => CLK_I, Q => 
                           n_2971, QN => n2686);
   KEY_EXPAN0_reg_21_24_inst : FD1 port map( D => n6162, CP => CLK_I, Q => 
                           n_2972, QN => n2689);
   KEY_EXPAN0_reg_20_24_inst : FD1 port map( D => n6161, CP => CLK_I, Q => 
                           n_2973, QN => n2688);
   KEY_EXPAN0_reg_19_24_inst : FD1 port map( D => n6160, CP => CLK_I, Q => 
                           n_2974, QN => n2691);
   KEY_EXPAN0_reg_18_24_inst : FD1 port map( D => n6159, CP => CLK_I, Q => 
                           n_2975, QN => n2690);
   KEY_EXPAN0_reg_17_24_inst : FD1 port map( D => n6158, CP => CLK_I, Q => 
                           n_2976, QN => n2693);
   KEY_EXPAN0_reg_16_24_inst : FD1 port map( D => n6157, CP => CLK_I, Q => 
                           n_2977, QN => n2692);
   KEY_EXPAN0_reg_15_24_inst : FD1 port map( D => n6156, CP => CLK_I, Q => 
                           n_2978, QN => n2679);
   KEY_EXPAN0_reg_14_24_inst : FD1 port map( D => n6155, CP => CLK_I, Q => 
                           n_2979, QN => n2678);
   KEY_EXPAN0_reg_13_24_inst : FD1 port map( D => n6154, CP => CLK_I, Q => 
                           n_2980, QN => n2681);
   KEY_EXPAN0_reg_12_24_inst : FD1 port map( D => n6153, CP => CLK_I, Q => 
                           n_2981, QN => n2680);
   KEY_EXPAN0_reg_11_24_inst : FD1 port map( D => n6152, CP => CLK_I, Q => 
                           n_2982, QN => n2683);
   KEY_EXPAN0_reg_10_24_inst : FD1 port map( D => n6151, CP => CLK_I, Q => 
                           n_2983, QN => n2682);
   KEY_EXPAN0_reg_9_24_inst : FD1 port map( D => n6150, CP => CLK_I, Q => 
                           n_2984, QN => n2685);
   KEY_EXPAN0_reg_8_24_inst : FD1 port map( D => n6149, CP => CLK_I, Q => 
                           n_2985, QN => n2684);
   KEY_EXPAN0_reg_7_24_inst : FD1 port map( D => n6148, CP => CLK_I, Q => 
                           n_2986, QN => n2671);
   KEY_EXPAN0_reg_6_24_inst : FD1 port map( D => n6147, CP => CLK_I, Q => 
                           n_2987, QN => n2670);
   KEY_EXPAN0_reg_5_24_inst : FD1 port map( D => n6146, CP => CLK_I, Q => 
                           n_2988, QN => n2673);
   KEY_EXPAN0_reg_4_24_inst : FD1 port map( D => n6145, CP => CLK_I, Q => 
                           n_2989, QN => n2672);
   KEY_EXPAN0_reg_3_24_inst : FD1 port map( D => n6144, CP => CLK_I, Q => 
                           n_2990, QN => n2675);
   KEY_EXPAN0_reg_2_24_inst : FD1 port map( D => n6143, CP => CLK_I, Q => 
                           n_2991, QN => n2674);
   KEY_EXPAN0_reg_1_24_inst : FD1 port map( D => n6142, CP => CLK_I, Q => 
                           n_2992, QN => n2677);
   KEY_EXPAN0_reg_0_24_inst : FD1 port map( D => n6141, CP => CLK_I, Q => 
                           n_2993, QN => n2676);
   v_KEY_COL_OUT0_reg_24_inst : FD1 port map( D => n4566, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_24_port, QN => n1867);
   v_TEMP_VECTOR_reg_16_inst : FD1 port map( D => n6693, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_16_port, QN => n_2994);
   KEY_EXPAN0_reg_63_16_inst : FD1 port map( D => n5692, CP => CLK_I, Q => 
                           n_2995, QN => n2599);
   KEY_EXPAN0_reg_62_16_inst : FD1 port map( D => n5691, CP => CLK_I, Q => 
                           n_2996, QN => n2598);
   KEY_EXPAN0_reg_61_16_inst : FD1 port map( D => n5690, CP => CLK_I, Q => 
                           n_2997, QN => n2601);
   KEY_EXPAN0_reg_60_16_inst : FD1 port map( D => n5689, CP => CLK_I, Q => 
                           n_2998, QN => n2600);
   KEY_EXPAN0_reg_59_16_inst : FD1 port map( D => n5688, CP => CLK_I, Q => 
                           n_2999, QN => n2603);
   KEY_EXPAN0_reg_58_16_inst : FD1 port map( D => n5687, CP => CLK_I, Q => 
                           n_3000, QN => n2602);
   KEY_EXPAN0_reg_57_16_inst : FD1 port map( D => n5686, CP => CLK_I, Q => 
                           n_3001, QN => n2605);
   KEY_EXPAN0_reg_56_16_inst : FD1 port map( D => n5685, CP => CLK_I, Q => 
                           n_3002, QN => n2604);
   KEY_EXPAN0_reg_55_16_inst : FD1 port map( D => n5684, CP => CLK_I, Q => 
                           n_3003, QN => n2591);
   KEY_EXPAN0_reg_54_16_inst : FD1 port map( D => n5683, CP => CLK_I, Q => 
                           n_3004, QN => n2590);
   KEY_EXPAN0_reg_53_16_inst : FD1 port map( D => n5682, CP => CLK_I, Q => 
                           n_3005, QN => n2593);
   KEY_EXPAN0_reg_52_16_inst : FD1 port map( D => n5681, CP => CLK_I, Q => 
                           n_3006, QN => n2592);
   KEY_EXPAN0_reg_51_16_inst : FD1 port map( D => n5680, CP => CLK_I, Q => 
                           n_3007, QN => n2595);
   KEY_EXPAN0_reg_50_16_inst : FD1 port map( D => n5679, CP => CLK_I, Q => 
                           n_3008, QN => n2594);
   KEY_EXPAN0_reg_49_16_inst : FD1 port map( D => n5678, CP => CLK_I, Q => 
                           n_3009, QN => n2597);
   KEY_EXPAN0_reg_48_16_inst : FD1 port map( D => n5677, CP => CLK_I, Q => 
                           n_3010, QN => n2596);
   KEY_EXPAN0_reg_47_16_inst : FD1 port map( D => n5676, CP => CLK_I, Q => 
                           n_3011, QN => n2583);
   KEY_EXPAN0_reg_46_16_inst : FD1 port map( D => n5675, CP => CLK_I, Q => 
                           n_3012, QN => n2582);
   KEY_EXPAN0_reg_45_16_inst : FD1 port map( D => n5674, CP => CLK_I, Q => 
                           n_3013, QN => n2585);
   KEY_EXPAN0_reg_44_16_inst : FD1 port map( D => n5673, CP => CLK_I, Q => 
                           n_3014, QN => n2584);
   KEY_EXPAN0_reg_43_16_inst : FD1 port map( D => n5672, CP => CLK_I, Q => 
                           n_3015, QN => n2587);
   KEY_EXPAN0_reg_42_16_inst : FD1 port map( D => n5671, CP => CLK_I, Q => 
                           n_3016, QN => n2586);
   KEY_EXPAN0_reg_41_16_inst : FD1 port map( D => n5670, CP => CLK_I, Q => 
                           n_3017, QN => n2589);
   KEY_EXPAN0_reg_40_16_inst : FD1 port map( D => n5669, CP => CLK_I, Q => 
                           n_3018, QN => n2588);
   KEY_EXPAN0_reg_39_16_inst : FD1 port map( D => n5668, CP => CLK_I, Q => 
                           n_3019, QN => n2575);
   KEY_EXPAN0_reg_38_16_inst : FD1 port map( D => n5667, CP => CLK_I, Q => 
                           n_3020, QN => n2574);
   KEY_EXPAN0_reg_37_16_inst : FD1 port map( D => n5666, CP => CLK_I, Q => 
                           n_3021, QN => n2577);
   KEY_EXPAN0_reg_36_16_inst : FD1 port map( D => n5665, CP => CLK_I, Q => 
                           n_3022, QN => n2576);
   KEY_EXPAN0_reg_35_16_inst : FD1 port map( D => n5664, CP => CLK_I, Q => 
                           n_3023, QN => n2579);
   KEY_EXPAN0_reg_34_16_inst : FD1 port map( D => n5663, CP => CLK_I, Q => 
                           n_3024, QN => n2578);
   KEY_EXPAN0_reg_33_16_inst : FD1 port map( D => n5662, CP => CLK_I, Q => 
                           n_3025, QN => n2581);
   KEY_EXPAN0_reg_32_16_inst : FD1 port map( D => n5661, CP => CLK_I, Q => 
                           n_3026, QN => n2580);
   KEY_EXPAN0_reg_31_16_inst : FD1 port map( D => n5660, CP => CLK_I, Q => 
                           n_3027, QN => n2631);
   KEY_EXPAN0_reg_30_16_inst : FD1 port map( D => n5659, CP => CLK_I, Q => 
                           n_3028, QN => n2630);
   KEY_EXPAN0_reg_29_16_inst : FD1 port map( D => n5658, CP => CLK_I, Q => 
                           n_3029, QN => n2633);
   KEY_EXPAN0_reg_28_16_inst : FD1 port map( D => n5657, CP => CLK_I, Q => 
                           n_3030, QN => n2632);
   KEY_EXPAN0_reg_27_16_inst : FD1 port map( D => n5656, CP => CLK_I, Q => 
                           n_3031, QN => n2635);
   KEY_EXPAN0_reg_26_16_inst : FD1 port map( D => n5655, CP => CLK_I, Q => 
                           n_3032, QN => n2634);
   KEY_EXPAN0_reg_25_16_inst : FD1 port map( D => n5654, CP => CLK_I, Q => 
                           n_3033, QN => n2637);
   KEY_EXPAN0_reg_24_16_inst : FD1 port map( D => n5653, CP => CLK_I, Q => 
                           n_3034, QN => n2636);
   KEY_EXPAN0_reg_23_16_inst : FD1 port map( D => n5652, CP => CLK_I, Q => 
                           n_3035, QN => n2623);
   KEY_EXPAN0_reg_22_16_inst : FD1 port map( D => n5651, CP => CLK_I, Q => 
                           n_3036, QN => n2622);
   KEY_EXPAN0_reg_21_16_inst : FD1 port map( D => n5650, CP => CLK_I, Q => 
                           n_3037, QN => n2625);
   KEY_EXPAN0_reg_20_16_inst : FD1 port map( D => n5649, CP => CLK_I, Q => 
                           n_3038, QN => n2624);
   KEY_EXPAN0_reg_19_16_inst : FD1 port map( D => n5648, CP => CLK_I, Q => 
                           n_3039, QN => n2627);
   KEY_EXPAN0_reg_18_16_inst : FD1 port map( D => n5647, CP => CLK_I, Q => 
                           n_3040, QN => n2626);
   KEY_EXPAN0_reg_17_16_inst : FD1 port map( D => n5646, CP => CLK_I, Q => 
                           n_3041, QN => n2629);
   KEY_EXPAN0_reg_16_16_inst : FD1 port map( D => n5645, CP => CLK_I, Q => 
                           n_3042, QN => n2628);
   KEY_EXPAN0_reg_15_16_inst : FD1 port map( D => n5644, CP => CLK_I, Q => 
                           n_3043, QN => n2615);
   KEY_EXPAN0_reg_14_16_inst : FD1 port map( D => n5643, CP => CLK_I, Q => 
                           n_3044, QN => n2614);
   KEY_EXPAN0_reg_13_16_inst : FD1 port map( D => n5642, CP => CLK_I, Q => 
                           n_3045, QN => n2617);
   KEY_EXPAN0_reg_12_16_inst : FD1 port map( D => n5641, CP => CLK_I, Q => 
                           n_3046, QN => n2616);
   KEY_EXPAN0_reg_11_16_inst : FD1 port map( D => n5640, CP => CLK_I, Q => 
                           n_3047, QN => n2619);
   KEY_EXPAN0_reg_10_16_inst : FD1 port map( D => n5639, CP => CLK_I, Q => 
                           n_3048, QN => n2618);
   KEY_EXPAN0_reg_9_16_inst : FD1 port map( D => n5638, CP => CLK_I, Q => 
                           n_3049, QN => n2621);
   KEY_EXPAN0_reg_8_16_inst : FD1 port map( D => n5637, CP => CLK_I, Q => 
                           n_3050, QN => n2620);
   KEY_EXPAN0_reg_7_16_inst : FD1 port map( D => n5636, CP => CLK_I, Q => 
                           n_3051, QN => n2607);
   KEY_EXPAN0_reg_6_16_inst : FD1 port map( D => n5635, CP => CLK_I, Q => 
                           n_3052, QN => n2606);
   KEY_EXPAN0_reg_5_16_inst : FD1 port map( D => n5634, CP => CLK_I, Q => 
                           n_3053, QN => n2609);
   KEY_EXPAN0_reg_4_16_inst : FD1 port map( D => n5633, CP => CLK_I, Q => 
                           n_3054, QN => n2608);
   KEY_EXPAN0_reg_3_16_inst : FD1 port map( D => n5632, CP => CLK_I, Q => 
                           n_3055, QN => n2611);
   KEY_EXPAN0_reg_2_16_inst : FD1 port map( D => n5631, CP => CLK_I, Q => 
                           n_3056, QN => n2610);
   KEY_EXPAN0_reg_1_16_inst : FD1 port map( D => n5630, CP => CLK_I, Q => 
                           n_3057, QN => n2613);
   KEY_EXPAN0_reg_0_16_inst : FD1 port map( D => n5629, CP => CLK_I, Q => 
                           n_3058, QN => n2612);
   v_KEY_COL_OUT0_reg_16_inst : FD1 port map( D => n4565, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_16_port, QN => n1929);
   v_TEMP_VECTOR_reg_8_inst : FD1 port map( D => n6701, CP => CLK_I, Q => 
                           v_TEMP_VECTOR_8_port, QN => n_3059);
   KEY_EXPAN0_reg_63_8_inst : FD1 port map( D => n5180, CP => CLK_I, Q => 
                           n_3060, QN => n2535);
   KEY_EXPAN0_reg_62_8_inst : FD1 port map( D => n5179, CP => CLK_I, Q => 
                           n_3061, QN => n2534);
   KEY_EXPAN0_reg_61_8_inst : FD1 port map( D => n5178, CP => CLK_I, Q => 
                           n_3062, QN => n2537);
   KEY_EXPAN0_reg_60_8_inst : FD1 port map( D => n5177, CP => CLK_I, Q => 
                           n_3063, QN => n2536);
   KEY_EXPAN0_reg_59_8_inst : FD1 port map( D => n5176, CP => CLK_I, Q => 
                           n_3064, QN => n2539);
   KEY_EXPAN0_reg_58_8_inst : FD1 port map( D => n5175, CP => CLK_I, Q => 
                           n_3065, QN => n2538);
   KEY_EXPAN0_reg_57_8_inst : FD1 port map( D => n5174, CP => CLK_I, Q => 
                           n_3066, QN => n2541);
   KEY_EXPAN0_reg_56_8_inst : FD1 port map( D => n5173, CP => CLK_I, Q => 
                           n_3067, QN => n2540);
   KEY_EXPAN0_reg_55_8_inst : FD1 port map( D => n5172, CP => CLK_I, Q => 
                           n_3068, QN => n2527);
   KEY_EXPAN0_reg_54_8_inst : FD1 port map( D => n5171, CP => CLK_I, Q => 
                           n_3069, QN => n2526);
   KEY_EXPAN0_reg_53_8_inst : FD1 port map( D => n5170, CP => CLK_I, Q => 
                           n_3070, QN => n2529);
   KEY_EXPAN0_reg_52_8_inst : FD1 port map( D => n5169, CP => CLK_I, Q => 
                           n_3071, QN => n2528);
   KEY_EXPAN0_reg_51_8_inst : FD1 port map( D => n5168, CP => CLK_I, Q => 
                           n_3072, QN => n2531);
   KEY_EXPAN0_reg_50_8_inst : FD1 port map( D => n5167, CP => CLK_I, Q => 
                           n_3073, QN => n2530);
   KEY_EXPAN0_reg_49_8_inst : FD1 port map( D => n5166, CP => CLK_I, Q => 
                           n_3074, QN => n2533);
   KEY_EXPAN0_reg_48_8_inst : FD1 port map( D => n5165, CP => CLK_I, Q => 
                           n_3075, QN => n2532);
   KEY_EXPAN0_reg_47_8_inst : FD1 port map( D => n5164, CP => CLK_I, Q => 
                           n_3076, QN => n2519);
   KEY_EXPAN0_reg_46_8_inst : FD1 port map( D => n5163, CP => CLK_I, Q => 
                           n_3077, QN => n2518);
   KEY_EXPAN0_reg_45_8_inst : FD1 port map( D => n5162, CP => CLK_I, Q => 
                           n_3078, QN => n2521);
   KEY_EXPAN0_reg_44_8_inst : FD1 port map( D => n5161, CP => CLK_I, Q => 
                           n_3079, QN => n2520);
   KEY_EXPAN0_reg_43_8_inst : FD1 port map( D => n5160, CP => CLK_I, Q => 
                           n_3080, QN => n2523);
   KEY_EXPAN0_reg_42_8_inst : FD1 port map( D => n5159, CP => CLK_I, Q => 
                           n_3081, QN => n2522);
   KEY_EXPAN0_reg_41_8_inst : FD1 port map( D => n5158, CP => CLK_I, Q => 
                           n_3082, QN => n2525);
   KEY_EXPAN0_reg_40_8_inst : FD1 port map( D => n5157, CP => CLK_I, Q => 
                           n_3083, QN => n2524);
   KEY_EXPAN0_reg_39_8_inst : FD1 port map( D => n5156, CP => CLK_I, Q => 
                           n_3084, QN => n2511);
   KEY_EXPAN0_reg_38_8_inst : FD1 port map( D => n5155, CP => CLK_I, Q => 
                           n_3085, QN => n2510);
   KEY_EXPAN0_reg_37_8_inst : FD1 port map( D => n5154, CP => CLK_I, Q => 
                           n_3086, QN => n2513);
   KEY_EXPAN0_reg_36_8_inst : FD1 port map( D => n5153, CP => CLK_I, Q => 
                           n_3087, QN => n2512);
   KEY_EXPAN0_reg_35_8_inst : FD1 port map( D => n5152, CP => CLK_I, Q => 
                           n_3088, QN => n2515);
   KEY_EXPAN0_reg_34_8_inst : FD1 port map( D => n5151, CP => CLK_I, Q => 
                           n_3089, QN => n2514);
   KEY_EXPAN0_reg_33_8_inst : FD1 port map( D => n5150, CP => CLK_I, Q => 
                           n_3090, QN => n2517);
   KEY_EXPAN0_reg_32_8_inst : FD1 port map( D => n5149, CP => CLK_I, Q => 
                           n_3091, QN => n2516);
   KEY_EXPAN0_reg_31_8_inst : FD1 port map( D => n5148, CP => CLK_I, Q => 
                           n_3092, QN => n2567);
   KEY_EXPAN0_reg_30_8_inst : FD1 port map( D => n5147, CP => CLK_I, Q => 
                           n_3093, QN => n2566);
   KEY_EXPAN0_reg_29_8_inst : FD1 port map( D => n5146, CP => CLK_I, Q => 
                           n_3094, QN => n2569);
   KEY_EXPAN0_reg_28_8_inst : FD1 port map( D => n5145, CP => CLK_I, Q => 
                           n_3095, QN => n2568);
   KEY_EXPAN0_reg_27_8_inst : FD1 port map( D => n5144, CP => CLK_I, Q => 
                           n_3096, QN => n2571);
   KEY_EXPAN0_reg_26_8_inst : FD1 port map( D => n5143, CP => CLK_I, Q => 
                           n_3097, QN => n2570);
   KEY_EXPAN0_reg_25_8_inst : FD1 port map( D => n5142, CP => CLK_I, Q => 
                           n_3098, QN => n2573);
   KEY_EXPAN0_reg_24_8_inst : FD1 port map( D => n5141, CP => CLK_I, Q => 
                           n_3099, QN => n2572);
   KEY_EXPAN0_reg_23_8_inst : FD1 port map( D => n5140, CP => CLK_I, Q => 
                           n_3100, QN => n2559);
   KEY_EXPAN0_reg_22_8_inst : FD1 port map( D => n5139, CP => CLK_I, Q => 
                           n_3101, QN => n2558);
   KEY_EXPAN0_reg_21_8_inst : FD1 port map( D => n5138, CP => CLK_I, Q => 
                           n_3102, QN => n2561);
   KEY_EXPAN0_reg_20_8_inst : FD1 port map( D => n5137, CP => CLK_I, Q => 
                           n_3103, QN => n2560);
   KEY_EXPAN0_reg_19_8_inst : FD1 port map( D => n5136, CP => CLK_I, Q => 
                           n_3104, QN => n2563);
   KEY_EXPAN0_reg_18_8_inst : FD1 port map( D => n5135, CP => CLK_I, Q => 
                           n_3105, QN => n2562);
   KEY_EXPAN0_reg_17_8_inst : FD1 port map( D => n5134, CP => CLK_I, Q => 
                           n_3106, QN => n2565);
   KEY_EXPAN0_reg_16_8_inst : FD1 port map( D => n5133, CP => CLK_I, Q => 
                           n_3107, QN => n2564);
   KEY_EXPAN0_reg_15_8_inst : FD1 port map( D => n5132, CP => CLK_I, Q => 
                           n_3108, QN => n2551);
   KEY_EXPAN0_reg_14_8_inst : FD1 port map( D => n5131, CP => CLK_I, Q => 
                           n_3109, QN => n2550);
   KEY_EXPAN0_reg_13_8_inst : FD1 port map( D => n5130, CP => CLK_I, Q => 
                           n_3110, QN => n2553);
   KEY_EXPAN0_reg_12_8_inst : FD1 port map( D => n5129, CP => CLK_I, Q => 
                           n_3111, QN => n2552);
   KEY_EXPAN0_reg_11_8_inst : FD1 port map( D => n5128, CP => CLK_I, Q => 
                           n_3112, QN => n2555);
   KEY_EXPAN0_reg_10_8_inst : FD1 port map( D => n5127, CP => CLK_I, Q => 
                           n_3113, QN => n2554);
   KEY_EXPAN0_reg_9_8_inst : FD1 port map( D => n5126, CP => CLK_I, Q => n_3114
                           , QN => n2557);
   KEY_EXPAN0_reg_8_8_inst : FD1 port map( D => n5125, CP => CLK_I, Q => n_3115
                           , QN => n2556);
   KEY_EXPAN0_reg_7_8_inst : FD1 port map( D => n5124, CP => CLK_I, Q => n_3116
                           , QN => n2543);
   KEY_EXPAN0_reg_6_8_inst : FD1 port map( D => n5123, CP => CLK_I, Q => n_3117
                           , QN => n2542);
   KEY_EXPAN0_reg_5_8_inst : FD1 port map( D => n5122, CP => CLK_I, Q => n_3118
                           , QN => n2545);
   KEY_EXPAN0_reg_4_8_inst : FD1 port map( D => n5121, CP => CLK_I, Q => n_3119
                           , QN => n2544);
   KEY_EXPAN0_reg_3_8_inst : FD1 port map( D => n5120, CP => CLK_I, Q => n_3120
                           , QN => n2547);
   KEY_EXPAN0_reg_2_8_inst : FD1 port map( D => n5119, CP => CLK_I, Q => n_3121
                           , QN => n2546);
   KEY_EXPAN0_reg_1_8_inst : FD1 port map( D => n5118, CP => CLK_I, Q => n_3122
                           , QN => n2549);
   KEY_EXPAN0_reg_0_8_inst : FD1 port map( D => n5117, CP => CLK_I, Q => n_3123
                           , QN => n2548);
   v_KEY_COL_OUT0_reg_8_inst : FD1 port map( D => n4564, CP => CLK_I, Q => 
                           v_KEY_COL_OUT0_8_port, QN => n1947);
   U149 : OR3 port map( A => n155, B => n156, C => n157, Z => n66);
   U161 : OR3 port map( A => n6676, B => n6675, C => n1833, Z => n179);
   U207 : OR2 port map( A => n6673, B => RESET_I, Z => n56);
   U267 : OR3 port map( A => n6792, B => n2391, C => n2091, Z => n275);
   U1896 : OR3 port map( A => n1587, B => n1873, C => n1874, Z => n1871);
   U1915 : AN3 port map( A => n2310, B => n6764, C => n1859, Z => n1926);
   U1917 : AN3 port map( A => n6740, B => n1932, C => n1933, Z => n1911);
   U1947 : AN3 port map( A => n2317, B => n1889, C => n6754, Z => n1997);
   U1982 : OR3 port map( A => n2308, B => n2321, C => n2039, Z => n2046);
   U1983 : OR2 port map( A => n6774, B => n2048, Z => n2045);
   U1984 : OR2 port map( A => n1843, B => n1977, Z => n2036);
   U2011 : OR2 port map( A => n2081, B => n2321, Z => n2078);
   U2033 : OR3 port map( A => n1897, B => n1763, C => n1936, Z => n2107);
   U2075 : AN3 port map( A => n2319, B => n6754, C => n1890, Z => n2159);
   U2120 : AN3 port map( A => n2201, B => n2202, C => n2203, Z => n2190);
   U2138 : AN3 port map( A => n2310, B => n6733, C => n1859, Z => n2221);
   U2145 : OR3 port map( A => n2111, B => n2314, C => n6776, Z => n2222);
   U2146 : OR3 port map( A => n2320, B => n2065, C => n2225, Z => n2213);
   U2250 : AN3 port map( A => n2319, B => n1903, C => n6733, Z => n2272);
   U2274 : AN3 port map( A => n2316, B => n2093, C => n1587, Z => n2278);
   U2362 : AN3 port map( A => n2301, B => n1877, C => n267, Z => n174);
   U2364 : AN3 port map( A => n1883, B => n1844, C => n2306, Z => n2301);
   U4512 : AN3 port map( A => n6654, B => n6655, C => n2487, Z => n2486);
   U4537 : AN3 port map( A => n6654, B => i_SRAM_ADDR_WR02, C => n2487, Z => 
                           n2488);
   U4562 : AN3 port map( A => n6655, B => i_SRAM_ADDR_WR01, C => n2487, Z => 
                           n2489);
   U4566 : AN3 port map( A => n6657, B => n6658, C => n6656, Z => n2470);
   U4570 : AN3 port map( A => n6657, B => i_SRAM_ADDR_WR05, C => n6656, Z => 
                           n2472);
   U4574 : AN3 port map( A => n6658, B => i_SRAM_ADDR_WR04, C => n6656, Z => 
                           n2473);
   U4578 : AN3 port map( A => i_SRAM_ADDR_WR05, B => i_SRAM_ADDR_WR04, C => 
                           n6656, Z => n2474);
   U4596 : AN4 port map( A => n2302, B => n6787, C => n2495, D => n2496, Z => 
                           n2493);
   U4600 : OR3 port map( A => n2299, B => v_CALCULATION_CNTR_2_port, C => n230,
                           Z => n2495);
   U4612 : AN3 port map( A => i_SRAM_ADDR_WR02, B => i_SRAM_ADDR_WR01, C => 
                           n2487, Z => n2490);
   U4635 : AN3 port map( A => n2306, B => n1883, C => v_CALCULATION_CNTR_4_port
                           , Z => n2498);
   U7 : NR2I port map( A => v_TEMP_VECTOR_31_port, B => n21, Z => n19);
   U12 : NR2I port map( A => v_TEMP_VECTOR_30_port, B => n21, Z => n26);
   U17 : NR2I port map( A => v_TEMP_VECTOR_29_port, B => n21, Z => n31);
   U22 : NR2I port map( A => v_TEMP_VECTOR_28_port, B => n21, Z => n36);
   U27 : NR2I port map( A => v_TEMP_VECTOR_27_port, B => n21, Z => n41);
   U32 : NR2I port map( A => v_TEMP_VECTOR_26_port, B => n21, Z => n46);
   U37 : NR2I port map( A => v_TEMP_VECTOR_25_port, B => n21, Z => n51);
   U40 : NR2I port map( A => n56, B => n57, Z => n18);
   U41 : NR2I port map( A => n1904, B => n2504, Z => n17);
   U45 : NR2I port map( A => v_TEMP_VECTOR_24_port, B => n21, Z => n60);
   U48 : ND2I port map( A => n64, B => n62, Z => n13);
   U49 : NR2I port map( A => n57, B => n65, Z => n64);
   U52 : ND2I port map( A => n6794, B => n2255, Z => n70);
   U57 : NR2I port map( A => v_TEMP_VECTOR_23_port, B => n80, Z => n78);
   U62 : NR2I port map( A => v_TEMP_VECTOR_22_port, B => n80, Z => n84);
   U67 : NR2I port map( A => v_TEMP_VECTOR_21_port, B => n80, Z => n88);
   U72 : NR2I port map( A => v_TEMP_VECTOR_20_port, B => n80, Z => n92);
   U77 : NR2I port map( A => v_TEMP_VECTOR_19_port, B => n80, Z => n96);
   U82 : NR2I port map( A => v_TEMP_VECTOR_18_port, B => n80, Z => n100);
   U87 : NR2I port map( A => v_TEMP_VECTOR_17_port, B => n80, Z => n104);
   U90 : NR2I port map( A => n108, B => n56, Z => n77);
   U91 : NR2I port map( A => n6784, B => n1904, Z => n76);
   U95 : NR2I port map( A => v_TEMP_VECTOR_16_port, B => n80, Z => n110);
   U98 : ND2I port map( A => n113, B => n112, Z => n73);
   U99 : NR2I port map( A => n108, B => n65, Z => n113);
   U105 : NR2I port map( A => v_TEMP_VECTOR_15_port, B => n121, Z => n119);
   U110 : NR2I port map( A => v_TEMP_VECTOR_14_port, B => n121, Z => n125);
   U115 : NR2I port map( A => v_TEMP_VECTOR_13_port, B => n121, Z => n129);
   U120 : NR2I port map( A => v_TEMP_VECTOR_12_port, B => n121, Z => n133);
   U125 : NR2I port map( A => v_TEMP_VECTOR_11_port, B => n121, Z => n137);
   U130 : NR2I port map( A => v_TEMP_VECTOR_10_port, B => n121, Z => n141);
   U135 : NR2I port map( A => v_TEMP_VECTOR_9_port, B => n121, Z => n145);
   U138 : NR2I port map( A => n149, B => n56, Z => n118);
   U139 : NR2I port map( A => n6782, B => n1904, Z => n117);
   U143 : NR2I port map( A => v_TEMP_VECTOR_8_port, B => n121, Z => n151);
   --U146 : NR2I port map( A => n154, B => n153, Z => n114);--changing NR2I with ND2I
   U146 : ND2I port map( A => n154, B => n153, Z => n114);
   U147 : NR2I port map( A => n149, B => n65, Z => n154);
   U152 : ND2I port map( A => n164, B => n165, Z => n160);
   U154 : ENI port map( A => v_KEY_COL_OUT0_7_port, B => v_TEMP_VECTOR_7_port, 
                           Z => n167);
   U155 : ENI port map( A => n169, B => v_TEMP_VECTOR_15_port, Z => n158);
   U160 : ENI port map( A => v_TEMP_VECTOR_14_port, B => n179, Z => n178);
   U162 : ENI port map( A => n2121, B => v_KEY_COL_OUT0_6_port, Z => n177);
   U166 : ND2I port map( A => n164, B => n184, Z => n182);
   U168 : ENI port map( A => v_KEY_COL_OUT0_5_port, B => v_TEMP_VECTOR_5_port, 
                           Z => n185);
   U169 : ENI port map( A => n186, B => v_TEMP_VECTOR_13_port, Z => n181);
   U173 : ND2I port map( A => n164, B => n191, Z => n189);
   U175 : ENI port map( A => v_KEY_COL_OUT0_4_port, B => v_TEMP_VECTOR_4_port, 
                           Z => n192);
   U177 : ENI port map( A => v_TEMP_VECTOR_12_port, B => n193, Z => n188);
   U181 : ND2I port map( A => n164, B => n197, Z => n195);
   U183 : ENI port map( A => v_KEY_COL_OUT0_3_port, B => v_TEMP_VECTOR_3_port, 
                           Z => n198);
   U184 : EOI port map( A => v_TEMP_VECTOR_11_port, B => n199, Z => n194);
   U188 : ND2I port map( A => n164, B => n205, Z => n203);
   U190 : ENI port map( A => v_KEY_COL_OUT0_2_port, B => v_TEMP_VECTOR_2_port, 
                           Z => n206);
   U191 : ENI port map( A => v_TEMP_VECTOR_10_port, B => n207, Z => n202);
   U193 : ND2I port map( A => n6675, B => n1875, Z => n208);
   U196 : ND2I port map( A => n164, B => n213, Z => n211);
   U198 : ND2I port map( A => n2304, B => n1904, Z => n168);
   U199 : ENI port map( A => v_KEY_COL_OUT0_1_port, B => v_TEMP_VECTOR_1_port, 
                           Z => n214);
   U200 : ENI port map( A => v_TEMP_VECTOR_9_port, B => n215, Z => n210);
   U201 : ND2I port map( A => n6674, B => n216, Z => n215);
   --U203 : AN2I port map( A => n164, B => n2325, Z => n159);-- changing AN2I with ND2I
   U203 : ND2I port map( A => n164, B => n2325, Z => n159);
   U206 : NR2I port map( A => n56, B => n6785, Z => n162);
   U210 : EOI port map( A => v_TEMP_VECTOR_8_port, B => n223, Z => n222);
   U213 : ENI port map( A => n2103, B => v_KEY_COL_OUT0_0_port, Z => n221);
   U214 : NR2I port map( A => n2325, B => n225, Z => n176);
   U215 : NR2I port map( A => n65, B => n6785, Z => n164);
   U233 : ND2I port map( A => n239, B => n231, Z => n233);
   U235 : ND2I port map( A => n240, B => n6802, Z => n231);
   U239 : ND2I port map( A => n1832, B => n1719, Z => n247);
   U241 : ND2I port map( A => n6789, B => n1877, Z => n252);
   U253 : ND2I port map( A => n239, B => n254, Z => n256);
   U259 : NR2I port map( A => n6786, B => n266, Z => n63);
   U262 : ND2I port map( A => n268, B => n6806, Z => n271);
   U264 : ND2I port map( A => n2479, B => n6806, Z => n273);
   U266 : ND2I port map( A => n274, B => n275, Z => n268);
   U269 : ND2I port map( A => n277, B => n6806, Z => n278);
   U271 : ND2I port map( A => n274, B => n280, Z => n277);
   U275 : NR2I port map( A => n4563, B => VALID_KEY_I, Z => n279);
   U279 : ND2I port map( A => n6676, B => n2050, Z => n187);
   U282 : ND2I port map( A => n6676, B => n1833, Z => n285);
   U287 : ND2I port map( A => n6674, B => n169, Z => n289);
   U289 : NR2I port map( A => n287, B => n65, Z => n282);
   U292 : ND2I port map( A => n6790, B => n2391, Z => n67);
   U333 : ND2I port map( A => n312, B => n2506, Z => n304);
   U351 : ND2I port map( A => n312, B => n2505, Z => n315);
   U372 : ND2I port map( A => n263, B => n1719, Z => n334);
   U376 : NR2I port map( A => n337, B => n338, Z => n336);
   U420 : NR2I port map( A => n445, B => n446, Z => n444);
   U464 : NR2I port map( A => n489, B => n490, Z => n488);
   U508 : NR2I port map( A => n533, B => n534, Z => n532);
   U552 : NR2I port map( A => n577, B => n578, Z => n576);
   U596 : NR2I port map( A => n621, B => n622, Z => n620);
   U640 : NR2I port map( A => n665, B => n666, Z => n664);
   U684 : NR2I port map( A => n709, B => n710, Z => n708);
   U728 : NR2I port map( A => n753, B => n754, Z => n752);
   U772 : NR2I port map( A => n797, B => n798, Z => n796);
   U816 : NR2I port map( A => n841, B => n842, Z => n840);
   U860 : NR2I port map( A => n885, B => n886, Z => n884);
   U904 : NR2I port map( A => n929, B => n930, Z => n928);
   U948 : NR2I port map( A => n973, B => n974, Z => n972);
   U992 : NR2I port map( A => n1017, B => n1018, Z => n1016);
   U1036 : NR2I port map( A => n1061, B => n1062, Z => n1060);
   U1080 : NR2I port map( A => n1105, B => n1106, Z => n1104);
   U1124 : NR2I port map( A => n1149, B => n1150, Z => n1148);
   U1168 : NR2I port map( A => n1193, B => n1194, Z => n1192);
   U1212 : NR2I port map( A => n1237, B => n1238, Z => n1236);
   U1256 : NR2I port map( A => n1281, B => n1282, Z => n1280);
   U1300 : NR2I port map( A => n1325, B => n1326, Z => n1324);
   U1344 : NR2I port map( A => n1369, B => n1370, Z => n1368);
   U1388 : NR2I port map( A => n1413, B => n1414, Z => n1412);
   U1432 : NR2I port map( A => n1457, B => n1458, Z => n1456);
   U1476 : NR2I port map( A => n1501, B => n1502, Z => n1500);
   U1520 : NR2I port map( A => n1545, B => n1546, Z => n1544);
   U1564 : NR2I port map( A => n1589, B => n1590, Z => n1588);
   U1608 : NR2I port map( A => n1633, B => n1634, Z => n1632);
   U1652 : NR2I port map( A => n1677, B => n1678, Z => n1676);
   U1696 : NR2I port map( A => n1721, B => n1722, Z => n1720);
   U1740 : NR2I port map( A => n1765, B => n1766, Z => n1764);
   U1749 : AN2I port map( A => n1780, B => n1781, Z => n1775);
   U1756 : AN2I port map( A => n1780, B => n1783, Z => n1782);
   U1764 : AN2I port map( A => n1780, B => n1789, Z => n1788);
   U1771 : AN2I port map( A => n1780, B => n1791, Z => n1790);
   U1772 : NR2I port map( A => n6801, B => n6800, Z => n1780);
   U1780 : AN2I port map( A => n1799, B => n1781, Z => n1798);
   U1787 : AN2I port map( A => n1799, B => n1783, Z => n1800);
   U1795 : AN2I port map( A => n1799, B => n1789, Z => n1805);
   U1802 : AN2I port map( A => n1799, B => n1791, Z => n1806);
   U1803 : NR2I port map( A => n1807, B => n6801, Z => n1799);
   U1813 : AN2I port map( A => n1781, B => n1818, Z => n1817);
   U1820 : AN2I port map( A => n1783, B => n1818, Z => n1819);
   U1828 : AN2I port map( A => n1789, B => n1818, Z => n1824);
   U1835 : AN2I port map( A => n1791, B => n1818, Z => n1825);
   U1836 : NR2I port map( A => n1808, B => n6800, Z => n1818);
   U1845 : AN2I port map( A => n1831, B => n1781, Z => n1830);
   --U1846 : AN2I port map( A => n6798, B => n6799, Z => n1781);--changing AN2I with NR2I
   U1846 : NR2I port map( A => n6798, B => n6799, Z => n1781);
   U1853 : AN2I port map( A => n1831, B => n1783, Z => n1834);
   U1854 : NR2I port map( A => n1835, B => n6799, Z => n1783);
   U1863 : AN2I port map( A => n1831, B => n1789, Z => n1841);
   U1864 : NR2I port map( A => n1836, B => n6798, Z => n1789);
   U1868 : NR2I port map( A => n6797, B => n6796, Z => n1776);
   U1870 : NR2I port map( A => n1845, B => n6797, Z => n1777);
   U1874 : NR2I port map( A => n1846, B => n6796, Z => n1778);
   U1877 : NR2I port map( A => n1845, B => n1846, Z => n1779);
   U1880 : AN2I port map( A => n1831, B => n1791, Z => n1842);
   U1881 : NR2I port map( A => n1836, B => n1835, Z => n1791);
   U1884 : NR2I port map( A => n1807, B => n1808, Z => n1831);
   U1889 : AO1P port map( A => n1849, B => n1850, C => n1851, D => n1852, Z => 
                      n1848);
   U1892 : ND2I port map( A => n6764, B => n6747, Z => n1860);
   U1893 : AN2I port map( A => n1863, B => n1864, Z => n1857);
   U1897 : ND2I port map( A => n6733, B => n1903, Z => n1869);
   U1906 : AO1P port map( A => n1763, B => n6746, C => n6767, D => n1907, Z => 
                           n1896);
   U1907 : NR2I port map( A => n6771, B => n6747, Z => n1907);
   U1911 : ND2I port map( A => n1901, B => n1918, Z => n1912);
   U1914 : AO1P port map( A => n1924, B => n6765, C => n1925, D => n1926, Z => 
                           n1919);
   U1928 : ND2I port map( A => n1959, B => n2320, Z => n1958);
   U1931 : ND2I port map( A => n6749, B => n6766, Z => n1965);
   U1940 : ND2I port map( A => n1985, B => n6766, Z => n1972);
   U1941 : AO1P port map( A => n1986, B => n2310, C => n1987, D => n1988, Z => 
                           n1955);
   U1943 : NR2I port map( A => n1887, B => n2321, Z => n1986);
   U1946 : AO1P port map( A => n2318, B => n1996, C => n1901, D => n1997, Z => 
                           n1995);
   U1948 : ND2I port map( A => n6671, B => n6730, Z => n1996);
   U1952 : AO1P port map( A => n2312, B => n1928, C => n2004, D => n2005, Z => 
                           n1990);
   U1956 : ND2I port map( A => n6764, B => n1864, Z => n1948);
   U1958 : NR2I port map( A => n2011, B => n1975, Z => n2007);
   U1961 : AO1P port map( A => n2013, B => n2014, C => n2015, D => n2016, Z => 
                           n2012);
   U1975 : ND2I port map( A => n6733, B => n6765, Z => n1928);
   U1989 : AO1P port map( A => n2310, B => n6730, C => n2056, D => n2057, Z => 
                           n2052);
   U1992 : AO1P port map( A => n1998, B => n6758, C => n2059, D => n2060, Z => 
                           n2014);
   U1994 : NR2I port map( A => n2063, B => n2048, Z => n2062);
   U1995 : NR2I port map( A => n1886, B => n1900, Z => n2061);
   U2004 : ND2I port map( A => n1850, B => n2320, Z => n2072);
   U2005 : AO1P port map( A => n2312, B => n2073, C => n2074, D => n2075, Z => 
                           n2071);
   U2013 : NR2I port map( A => n1850, B => n1901, Z => n2026);
   U2019 : ND2I port map( A => n1859, B => n2093, Z => n2092);
   U2026 : ND2I port map( A => n1909, B => n1763, Z => n2104);
   U2028 : ND2I port map( A => n2105, B => n2305, Z => n1870);
   U2035 : AO1P port map( A => n1915, B => n2312, C => n2112, D => n2113, Z => 
                           n2094);
   U2037 : ND2I port map( A => n2116, B => n2117, Z => n2112);
   U2043 : ND2I port map( A => n4561, B => n2391, Z => n2123);
   U2048 : ND2I port map( A => n2130, B => n2131, Z => n2126);
   U2051 : ND2I port map( A => n1970, B => n6760, Z => n1973);
   U2065 : AO1P port map( A => n2147, B => n1924, C => n2148, D => n2149, Z => 
                           n2145);
   U2072 : NR2I port map( A => n1587, B => n2305, Z => n2154);
   U2074 : AO1P port map( A => n2318, B => n6750, C => n2158, D => n2159, Z => 
                           n2157);
   U2076 : AN2I port map( A => n2315, B => n2147, Z => n2158);
   U2077 : NR2I port map( A => n2051, B => n2084, Z => n2147);
   U2081 : ND2I port map( A => n6764, B => n1903, Z => n2160);
   U2086 : AO1P port map( A => n1886, B => n1889, C => n2173, D => n2174, Z => 
                           n2172);
   U2088 : ND2I port map( A => n1763, B => n2308, Z => n2176);
   U2090 : ND2I port map( A => n1890, B => n6759, Z => n2073);
   U2093 : ND2I port map( A => n6747, B => n6759, Z => n2032);
   U2098 : ND2I port map( A => n1900, B => n2114, Z => n2179);
   U2099 : ND2I port map( A => n1874, B => n6757, Z => n2114);
   U2100 : NR2I port map( A => n2182, B => n2063, Z => n2054);
   U2105 : NR2I port map( A => n1889, B => n2025, Z => n2011);
   U2108 : NR2I port map( A => n6774, B => n1859, Z => n1988);
   U2109 : ND2I port map( A => n1953, B => n2189, Z => n2163);
   U2113 : ND2I port map( A => n1937, B => n1889, Z => n2196);
   U2121 : AO1P port map( A => n2204, B => n6770, C => n2206, D => n2207, Z => 
                           n2203);
   U2125 : ENI port map( A => n1858, B => n1897, Z => n2039);
   U2126 : NR2I port map( A => n6768, B => n6775, Z => n2204);
   U2129 : NR2I port map( A => n1887, B => n1944, Z => n1977);
   U2132 : ND2I port map( A => n1953, B => n2211, Z => n2210);
   U2137 : NR2I port map( A => n2151, B => n2221, Z => n2218);
   U2139 : NR2I port map( A => n1936, B => n6774, Z => n2151);
   U2142 : ND2I port map( A => n6671, B => n2224, Z => n2119);
   U2144 : NR2I port map( A => n2048, B => n1944, Z => n1895);
   U2150 : NR2I port map( A => n2316, B => n2084, Z => n2055);
   U2151 : NR2I port map( A => n2314, B => n1858, Z => n2084);
   U2155 : NR2I port map( A => n1897, B => n2311, Z => n2105);
   U2158 : NR2I port map( A => n2081, B => n6747, Z => n2228);
   U2160 : ND2I port map( A => n1970, B => n6749, Z => n2049);
   U2162 : NR2I port map( A => n1878, B => n1763, Z => n1886);
   U2168 : ND2I port map( A => n6764, B => n6757, Z => n2238);
   U2171 : NR2I port map( A => n6771, B => n1969, Z => n2141);
   U2174 : NR2I port map( A => n6774, B => n6772, Z => n1946);
   U2177 : ND2I port map( A => n1864, B => n1985, Z => n2118);
   U2180 : ND2I port map( A => n1936, B => n6671, Z => n2003);
   U2181 : AO1P port map( A => n2319, B => n2155, C => n2242, D => n2243, Z => 
                           n2229);
   U2183 : ND2I port map( A => n1763, B => n6750, Z => n2245);
   U2187 : ND2I port map( A => n1874, B => n6766, Z => n2155);
   U2189 : NR2I port map( A => n2025, B => n6768, Z => n2000);
   U2192 : ND2I port map( A => n1951, B => n2250, Z => n2249);
   U2197 : NR2I port map( A => n1938, B => n2198, Z => n1915);
   U2198 : ND2I port map( A => n6671, B => n2106, Z => n2115);
   U2199 : ND2I port map( A => n2314, B => n1858, Z => n2106);
   U2201 : NR2I port map( A => n1858, B => n6755, Z => n2182);
   U2204 : NR2I port map( A => n2187, B => n2063, Z => n2178);
   U2205 : NR2I port map( A => n1885, B => n2025, Z => n2063);
   U2208 : ND2I port map( A => n1864, B => n6744, Z => n2077);
   U2210 : NR2I port map( A => n2208, B => n2198, Z => n1909);
   U2212 : ND2I port map( A => n1874, B => n6739, Z => n2129);
   U2213 : ND2I port map( A => n2314, B => n2025, Z => n1874);
   U2214 : NR2I port map( A => n1938, B => n1944, Z => n1894);
   U2215 : NR2I port map( A => n2305, B => n2314, Z => n1944);
   U2216 : NR2I port map( A => n2320, B => n1873, Z => n1980);
   U2222 : ND2I port map( A => n1970, B => n1985, Z => n2140);
   U2223 : ND2I port map( A => n2316, B => n2025, Z => n1985);
   U2224 : ND2I port map( A => n1858, B => n6751, Z => n1970);
   U2227 : ND2I port map( A => n6765, B => n6749, Z => n2241);
   U2229 : NR2I port map( A => n6751, B => n1858, Z => n2188);
   U2231 : ND2I port map( A => n2024, B => n6768, Z => n2102);
   U2234 : NR2I port map( A => n2305, B => n2321, Z => n2051);
   U2235 : NR2I port map( A => n1890, B => n1858, Z => n2187);
   U2237 : ND2I port map( A => n1998, B => n1936, Z => n2264);
   U2238 : ND2I port map( A => n6755, B => n1858, Z => n1936);
   U2239 : ND2I port map( A => n2313, B => n2093, Z => n1898);
   U2240 : NR2I port map( A => n2391, B => n4558, Z => n1951);
   U2243 : ND2I port map( A => n1901, B => n2269, Z => n2268);
   U2245 : AO1P port map( A => n2318, B => n6755, C => n2272, D => n2273, Z => 
                           n2271);
   U2249 : NR2I port map( A => n2197, B => n1858, Z => n1887);
   U2253 : NR2I port map( A => n6776, B => n1763, Z => n1902);
   U2254 : NR2I port map( A => n1858, B => n2321, Z => n2111);
   U2255 : NR2I port map( A => n1969, B => n6768, Z => n1976);
   U2256 : ND2I port map( A => n6769, B => n6739, Z => n2090);
   U2258 : NR2I port map( A => n2025, B => n6747, Z => n1940);
   U2261 : ND2I port map( A => n6733, B => n2224, Z => n2058);
   U2263 : NR2I port map( A => n6779, B => n1878, Z => n1916);
   U2264 : NR2I port map( A => n2048, B => n2198, Z => n2246);
   U2265 : NR2I port map( A => n6751, B => n2305, Z => n2198);
   U2266 : NR2I port map( A => n6779, B => n6774, Z => n1914);
   U2268 : NR2I port map( A => n2320, B => n1763, Z => n2184);
   U2270 : ND2I port map( A => n6747, B => n1863, Z => n1930);
   U2271 : ND2I port map( A => n6751, B => n2025, Z => n1863);
   U2273 : AO1P port map( A => n2028, B => n1998, C => n1901, D => n2278, Z => 
                           n2277);
   U2276 : ND2I port map( A => n2279, B => n2280, Z => n1893);
   U2279 : NR2I port map( A => n6774, B => n1763, Z => n1998);
   U2280 : NR2I port map( A => n1938, B => n2083, Z => n2028);
   U2281 : NR2I port map( A => n2025, B => n2316, Z => n2083);
   U2282 : NR2I port map( A => n1885, B => n1858, Z => n1938);
   U2284 : NR2I port map( A => n6774, B => n2311, Z => n1881);
   U2286 : NR2I port map( A => n1897, B => n1587, Z => n1937);
   U2287 : NR2I port map( A => n6776, B => n2311, Z => n1945);
   U2289 : NR2I port map( A => n2308, B => n1897, Z => n1924);
   U2290 : NR2I port map( A => n6768, B => n1858, Z => n2048);
   U2292 : NR2I port map( A => n1675, B => n2311, Z => n1934);
   U2294 : ND2I port map( A => n6733, B => n1864, Z => n2239);
   U2295 : ND2I port map( A => n1858, B => n1969, Z => n1864);
   U2297 : NR2I port map( A => n1858, B => n2316, Z => n1975);
   U2298 : NR2I port map( A => n1885, B => n6755, Z => n2006);
   U2299 : NR2I port map( A => n2311, B => n1878, Z => n1900);
   U2303 : NR2I port map( A => n6772, B => n2314, Z => n2043);
   U2305 : NR2I port map( A => n2305, B => n1763, Z => n2024);
   U2306 : NR2I port map( A => n1763, B => n1858, Z => n2093);
   U2309 : NR2I port map( A => n1969, B => n1885, Z => n2020);
   U2311 : NR2I port map( A => n1587, B => n6777, Z => n2044);
   U2314 : NR2I port map( A => n1675, B => n1763, Z => n1923);
   U2316 : ND2I port map( A => n2283, B => n2284, Z => n1873);
   U2320 : NR2I port map( A => n2308, B => n6777, Z => n1927);
   U2325 : ND2I port map( A => n2287, B => n2288, Z => n2047);
   U2328 : ND2I port map( A => n6744, B => n2224, Z => n1983);
   U2329 : ND2I port map( A => n1858, B => n6747, Z => n2224);
   U2331 : NR2I port map( A => n6747, B => n1858, Z => n2208);
   U2333 : ND2I port map( A => n2289, B => n2290, Z => n2025);
   U2337 : NR2I port map( A => n6755, B => n6768, Z => n2197);
   U2339 : ND2I port map( A => n2291, B => n2292, Z => n1885);
   U2346 : NR2I port map( A => n1850, B => n2391, Z => n1953);
   U2347 : ND2I port map( A => n2295, B => n2296, Z => n1850);
   U2350 : ND2I port map( A => v_CALCULATION_CNTR_1_port, B => n2255, Z => 
                           n2298);
   U2353 : ND2I port map( A => n6794, B => n1882, Z => n2300);
   U2355 : ND2I port map( A => v_CALCULATION_CNTR_2_port, B => n2301, Z => n266
                           );
   U2358 : ND2I port map( A => n2302, B => n2303, Z => n2281);
   U2361 : NR2I port map( A => n225, B => n174, Z => n166);
   U2363 : NR2I port map( A => n2255, B => n1882, Z => n267);
   U2370 : NR2I port map( A => n6804, B => n2391, Z => n263);
   U4487 : ND2I port map( A => n6653, B => n2485, Z => n2480);
   U4598 : ND2I port map( A => n2498, B => n2299, Z => n68);
   U4599 : NR2I port map( A => v_CALCULATION_CNTR_2_port, B => n1882, Z => 
                           n2497);
   U4602 : ND2I port map( A => n2307, B => n2299, Z => n2302);
   U4603 : NR2I port map( A => v_CALCULATION_CNTR_1_port, B => 
                           v_CALCULATION_CNTR_0_port, Z => n2299);
   U4604 : NR2I port map( A => n230, B => n1877, Z => n2307);
   U4613 : NR2I port map( A => n6802, B => n6653, Z => n2487);
   U4615 : NR2I port map( A => n2391, B => n2509, Z => n2485);
   U4639 : ND2I port map( A => n6673, B => n6806, Z => n65);
   U4642 : ND2I port map( A => n2391, B => n6806, Z => n242);
   U4645 : NR2I port map( A => n1793, B => n1974, Z => KEY_EXP_O(9));
   U4647 : NR2I port map( A => n1793, B => n1947, Z => KEY_EXP_O(8));
   U4649 : NR2I port map( A => n1793, B => n1866, Z => KEY_EXP_O(7));
   U4651 : NR2I port map( A => n1793, B => n1861, Z => KEY_EXP_O(6));
   U4653 : NR2I port map( A => n1793, B => n1906, Z => KEY_EXP_O(5));
   U4655 : NR2I port map( A => n1793, B => n2023, Z => KEY_EXP_O(4));
   U4657 : NR2I port map( A => n1793, B => n2001, Z => KEY_EXP_O(3));
   U4659 : NR2I port map( A => n1793, B => n1941, Z => KEY_EXP_O(31));
   U4661 : NR2I port map( A => n1793, B => n1865, Z => KEY_EXP_O(30));
   U4663 : NR2I port map( A => n1793, B => n1968, Z => KEY_EXP_O(2));
   U4665 : NR2I port map( A => n1793, B => n1921, Z => KEY_EXP_O(29));
   U4667 : NR2I port map( A => n1793, B => n1967, Z => KEY_EXP_O(28));
   U4669 : NR2I port map( A => n1793, B => n1868, Z => KEY_EXP_O(27));
   U4671 : NR2I port map( A => n1793, B => n1999, Z => KEY_EXP_O(26));
   U4673 : NR2I port map( A => n1793, B => n1989, Z => KEY_EXP_O(25));
   U4675 : NR2I port map( A => n1793, B => n1867, Z => KEY_EXP_O(24));
   U4677 : NR2I port map( A => n1793, B => n1917, Z => KEY_EXP_O(23));
   U4679 : NR2I port map( A => n1793, B => n1910, Z => KEY_EXP_O(22));
   U4681 : NR2I port map( A => n1793, B => n1931, Z => KEY_EXP_O(21));
   U4683 : NR2I port map( A => n1793, B => n1984, Z => KEY_EXP_O(20));
   U4685 : NR2I port map( A => n1793, B => n1966, Z => KEY_EXP_O(1));
   U4687 : NR2I port map( A => n1793, B => n1962, Z => KEY_EXP_O(19));
   U4689 : NR2I port map( A => n1793, B => n1956, Z => KEY_EXP_O(18));
   U4691 : NR2I port map( A => n1793, B => n1949, Z => KEY_EXP_O(17));
   U4693 : NR2I port map( A => n1793, B => n1929, Z => KEY_EXP_O(16));
   U4695 : NR2I port map( A => n1793, B => n1908, Z => KEY_EXP_O(15));
   U4697 : NR2I port map( A => n1793, B => n1862, Z => KEY_EXP_O(14));
   U4699 : NR2I port map( A => n1793, B => n1905, Z => KEY_EXP_O(13));
   U4701 : NR2I port map( A => n1793, B => n1982, Z => KEY_EXP_O(12));
   U4703 : NR2I port map( A => n1793, B => n1872, Z => KEY_EXP_O(11));
   U4705 : NR2I port map( A => n1793, B => n1922, Z => KEY_EXP_O(10));
   U4707 : NR2I port map( A => n1793, B => n1981, Z => KEY_EXP_O(0));
   U3 : ND2I port map( A => n1805, B => n1777, Z => n1);
   U4 : ND2I port map( A => n1788, B => n1777, Z => n2);
   U5 : ND2I port map( A => n1775, B => n1777, Z => n3);
   U6 : ND2I port map( A => n1788, B => n1776, Z => n4);
   U8 : ND2I port map( A => n1775, B => n1776, Z => n5);
   U9 : ND2I port map( A => n1841, B => n1779, Z => n6);
   U10 : ND2I port map( A => n1830, B => n1779, Z => n7);
   U11 : ND2I port map( A => n1834, B => n1779, Z => n8);
   U13 : ND2I port map( A => n1817, B => n1779, Z => n9);
   U14 : ND2I port map( A => n1805, B => n1779, Z => n10);
   U15 : ND2I port map( A => n1798, B => n1779, Z => n11);
   U16 : ND2I port map( A => n1788, B => n1779, Z => n12);
   U18 : ND2I port map( A => n1824, B => n1778, Z => n14);
   U19 : ND2I port map( A => n1805, B => n1778, Z => n22);
   U20 : ND2I port map( A => n1788, B => n1778, Z => n23);
   U21 : ND2I port map( A => n1824, B => n1779, Z => n28);
   U23 : ND2I port map( A => n1798, B => n1776, Z => n33);
   U24 : ND2I port map( A => n1805, B => n1776, Z => n38);
   U25 : ND2I port map( A => n1798, B => n1777, Z => n43);
   U26 : ND2I port map( A => n1842, B => n1779, Z => n48);
   U28 : ND2I port map( A => n1825, B => n1779, Z => n53);
   U29 : ND2I port map( A => n1779, B => n1819, Z => n58);
   U30 : ND2I port map( A => n1806, B => n1779, Z => n59);
   U31 : ND2I port map( A => n1800, B => n1779, Z => n69);
   U33 : ND2I port map( A => n1790, B => n1779, Z => n71);
   U34 : ND2I port map( A => n1775, B => n1779, Z => n72);
   U35 : ND2I port map( A => n1782, B => n1779, Z => n81);
   U36 : ND2I port map( A => n1841, B => n1778, Z => n109);
   U38 : ND2I port map( A => n1842, B => n1778, Z => n122);
   U39 : ND2I port map( A => n1830, B => n1778, Z => n150);
   U42 : ND2I port map( A => n1834, B => n1778, Z => n163);
   U43 : ND2I port map( A => n1825, B => n1778, Z => n170);
   U44 : ND2I port map( A => n1817, B => n1778, Z => n180);
   U46 : ND2I port map( A => n1778, B => n1819, Z => n200);
   U47 : ND2I port map( A => n1806, B => n1778, Z => n209);
   U50 : ND2I port map( A => n1798, B => n1778, Z => n217);
   U51 : ND2I port map( A => n1800, B => n1778, Z => n224);
   U53 : ND2I port map( A => n1790, B => n1778, Z => n227);
   U54 : ND2I port map( A => n1775, B => n1778, Z => n228);
   U55 : ND2I port map( A => n1782, B => n1778, Z => n229);
   U56 : ND2I port map( A => n1841, B => n1777, Z => n232);
   U58 : ND2I port map( A => n1841, B => n1776, Z => n234);
   U59 : ND2I port map( A => n1830, B => n1777, Z => n235);
   U60 : ND2I port map( A => n1830, B => n1776, Z => n236);
   U61 : ND2I port map( A => n1824, B => n1777, Z => n237);
   U63 : ND2I port map( A => n1824, B => n1776, Z => n238);
   U64 : ND2I port map( A => n1817, B => n1777, Z => n241);
   U65 : ND2I port map( A => n1817, B => n1776, Z => n245);
   U66 : ND2I port map( A => n1842, B => n1777, Z => n246);
   U68 : ND2I port map( A => n1842, B => n1776, Z => n248);
   U69 : ND2I port map( A => n1825, B => n1777, Z => n249);
   U70 : ND2I port map( A => n1825, B => n1776, Z => n250);
   U71 : ND2I port map( A => n1806, B => n1777, Z => n251);
   U73 : ND2I port map( A => n1806, B => n1776, Z => n253);
   U74 : ND2I port map( A => n1790, B => n1777, Z => n255);
   U75 : ND2I port map( A => n1790, B => n1776, Z => n257);
   U76 : ND2I port map( A => n1834, B => n1777, Z => n258);
   U78 : ND2I port map( A => n1834, B => n1776, Z => n259);
   U79 : ND2I port map( A => n1777, B => n1819, Z => n260);
   U80 : ND2I port map( A => n1776, B => n1819, Z => n261);
   U81 : ND2I port map( A => n1800, B => n1777, Z => n265);
   U83 : ND2I port map( A => n1800, B => n1776, Z => n269);
   U84 : ND2I port map( A => n1782, B => n1777, Z => n270);
   U85 : ND2I port map( A => n1782, B => n1776, Z => n272);
   U86 : IVDA port map( A => n2469, Y => n_3124, Z => n276);
   U88 : IVDA port map( A => n2461, Y => n_3125, Z => n284);
   U89 : IVDA port map( A => n2468, Y => n_3126, Z => n286);
   U92 : IVDA port map( A => n2460, Y => n_3127, Z => n293);
   U93 : IVDA port map( A => n2467, Y => n_3128, Z => n301);
   U94 : IVDA port map( A => n2459, Y => n_3129, Z => n303);
   U96 : IVDA port map( A => n2466, Y => n_3130, Z => n314);
   U97 : IVDA port map( A => n2458, Y => n_3131, Z => n325);
   U100 : IVDA port map( A => n2465, Y => n_3132, Z => n335);
   U101 : IVDA port map( A => n2457, Y => n_3133, Z => n347);
   U102 : IVDA port map( A => n2464, Y => n_3134, Z => n348);
   U103 : IVDA port map( A => n2456, Y => n_3135, Z => n349);
   U104 : IVDA port map( A => n2463, Y => n_3136, Z => n350);
   U106 : IVDA port map( A => n2462, Y => n_3137, Z => n351);
   U107 : IVDA port map( A => n2440, Y => n_3138, Z => n352);
   U108 : IVDA port map( A => n2309, Y => n_3139, Z => n353);
   U109 : IVDA port map( A => n2445, Y => n_3140, Z => n354);
   U111 : IVDA port map( A => n2453, Y => n_3141, Z => n359);
   U112 : IVDA port map( A => n2444, Y => n_3142, Z => n360);
   U113 : IVDA port map( A => n2452, Y => n_3143, Z => n361);
   U114 : IVDA port map( A => n2443, Y => n_3144, Z => n362);
   U116 : IVDA port map( A => n2451, Y => n_3145, Z => n363);
   U117 : IVDA port map( A => n2442, Y => n_3146, Z => n364);
   U118 : IVDA port map( A => n2450, Y => n_3147, Z => n365);
   U119 : IVDA port map( A => n2449, Y => n_3148, Z => n366);
   U121 : IVDA port map( A => n2448, Y => n_3149, Z => n371);
   U122 : IVDA port map( A => n2455, Y => n_3150, Z => n372);
   U123 : IVDA port map( A => n2447, Y => n_3151, Z => n373);
   U124 : IVDA port map( A => n2454, Y => n_3152, Z => n374);
   U126 : IVDA port map( A => n2446, Y => n_3153, Z => n375);
   U127 : IVDA port map( A => n2441, Y => n_3154, Z => n376);
   U128 : IVDA port map( A => n2439, Y => n_3155, Z => n377);
   U129 : AO4 port map( A => n6657, B => n231, C => n2297, D => n233, Z => 
                           n6713);
   U131 : AO4 port map( A => n6663, B => n254, C => n2274, D => n256, Z => 
                           n6721);
   U132 : EON1 port map( A => n1882, B => n242, C => N1748, D => n2499, Z => 
                           n6666);
   U133 : AN2I port map( A => n2470, B => n2471, Z => n378);
   U134 : AN2I port map( A => n2472, B => n2471, Z => n383);
   U136 : AN2I port map( A => n2473, B => n2471, Z => n384);
   U137 : AN2I port map( A => n2474, B => n2471, Z => n385);
   U140 : AN2I port map( A => n2475, B => n2471, Z => n386);
   U141 : AN2I port map( A => n2476, B => n2471, Z => n387);
   U142 : AN2I port map( A => n2477, B => n2471, Z => n388);
   U144 : AN2I port map( A => n2478, B => n2471, Z => n389);
   U145 : AN2I port map( A => n2482, B => n2470, Z => n390);
   U148 : AN2I port map( A => n2482, B => n2472, Z => n399);
   U150 : AN2I port map( A => n2482, B => n2473, Z => n400);
   U151 : AN2I port map( A => n2482, B => n2474, Z => n401);
   U153 : AN2I port map( A => n2482, B => n2475, Z => n402);
   U156 : AN2I port map( A => n2482, B => n2476, Z => n403);
   U157 : AN2I port map( A => n2482, B => n2477, Z => n404);
   U158 : AN2I port map( A => n2482, B => n2478, Z => n405);
   U159 : AN2I port map( A => n2483, B => n2470, Z => n406);
   U163 : AN2I port map( A => n2483, B => n2472, Z => n411);
   U164 : AN2I port map( A => n2483, B => n2473, Z => n412);
   U165 : AN2I port map( A => n2483, B => n2474, Z => n413);
   U167 : AN2I port map( A => n2483, B => n2475, Z => n414);
   U170 : AN2I port map( A => n2483, B => n2476, Z => n415);
   U171 : AN2I port map( A => n2483, B => n2477, Z => n416);
   U172 : AN2I port map( A => n2483, B => n2478, Z => n417);
   U174 : AN2I port map( A => n2484, B => n2470, Z => n418);
   U176 : AN2I port map( A => n2484, B => n2472, Z => n423);
   U178 : AN2I port map( A => n2484, B => n2473, Z => n424);
   U179 : AN2I port map( A => n2484, B => n2474, Z => n425);
   U180 : AN2I port map( A => n2484, B => n2475, Z => n426);
   U182 : AN2I port map( A => n2484, B => n2476, Z => n427);
   U185 : AN2I port map( A => n2484, B => n2477, Z => n428);
   U186 : AN2I port map( A => n2484, B => n2478, Z => n429);
   U187 : AN2I port map( A => n2486, B => n2475, Z => n430);
   U189 : AN2I port map( A => n2486, B => n2476, Z => n435);
   U192 : AN2I port map( A => n2486, B => n2477, Z => n436);
   U194 : AN2I port map( A => n2486, B => n2478, Z => n437);
   U195 : AN2I port map( A => n2488, B => n2475, Z => n438);
   U197 : AN2I port map( A => n2488, B => n2476, Z => n439);
   U202 : AN2I port map( A => n2488, B => n2477, Z => n440);
   U204 : AN2I port map( A => n2488, B => n2478, Z => n441);
   U205 : AN2I port map( A => n2489, B => n2475, Z => n442);
   U208 : AN2I port map( A => n2489, B => n2476, Z => n443);
   U209 : AN2I port map( A => n2489, B => n2477, Z => n487);
   U211 : AN2I port map( A => n2489, B => n2478, Z => n531);
   U212 : AN2I port map( A => n2490, B => n2475, Z => n575);
   U216 : AN2I port map( A => n2490, B => n2476, Z => n619);
   U217 : AN2I port map( A => n2490, B => n2477, Z => n663);
   U218 : AN2I port map( A => n2490, B => n2478, Z => n707);
   U219 : AN2I port map( A => n2486, B => n2470, Z => n751);
   U220 : AN2I port map( A => n2486, B => n2472, Z => n795);
   U221 : AN2I port map( A => n2486, B => n2473, Z => n839);
   U222 : AN2I port map( A => n2486, B => n2474, Z => n883);
   U223 : AN2I port map( A => n2488, B => n2470, Z => n927);
   U224 : AN2I port map( A => n2488, B => n2472, Z => n971);
   U225 : AN2I port map( A => n2488, B => n2473, Z => n1015);
   U226 : AN2I port map( A => n2488, B => n2474, Z => n1059);
   U227 : AN2I port map( A => n2489, B => n2470, Z => n1103);
   U228 : AN2I port map( A => n2489, B => n2472, Z => n1147);
   U229 : AN2I port map( A => n2489, B => n2473, Z => n1191);
   U230 : AN2I port map( A => n2489, B => n2474, Z => n1235);
   U231 : AN2I port map( A => n2490, B => n2470, Z => n1279);
   U232 : AN2I port map( A => n2490, B => n2472, Z => n1323);
   U234 : AN2I port map( A => n2490, B => n2473, Z => n1367);
   U236 : AN2I port map( A => n2490, B => n2474, Z => n1411);
   U237 : NR2I port map( A => n1543, B => n2493, Z => n1499);
   U238 : NR3 port map( A => n1832, B => n4563, C => n1719, Z => n1543);
   U240 : NR2I port map( A => n2197, B => n2314, Z => n1859);
   U242 : ENI port map( A => i_INTERN_ADDR_RD0, B => n2395, Z => n2098);
   U243 : ENI port map( A => i_SRAM_ADDR_WR0, B => n2399, Z => n2101);
   U244 : EOI port map( A => i_INTERN_ADDR_RD01, B => n2394, Z => n2127);
   U245 : ENI port map( A => i_INTERN_ADDR_RD02, B => n2393, Z => n2134);
   U246 : EOI port map( A => i_SRAM_ADDR_WR01, B => n2398, Z => n2146);
   U247 : ENI port map( A => i_SRAM_ADDR_WR02, B => n2397, Z => n2150);
   U248 : EOI port map( A => i_INTERN_ADDR_RD03, B => n2392, Z => n2175);
   U249 : EOI port map( A => i_SRAM_ADDR_WR03, B => n2396, Z => n2177);
   U250 : AO4 port map( A => n1792, B => n1973, C => n6741, D => n1631, Z => 
                           n2087);
   U251 : AO4 port map( A => n1972, B => n6773, C => n1973, D => n6775, Z => 
                           n1971);
   U252 : AO2 port map( A => n1998, B => n6747, C => n1886, D => n6734, Z => 
                           n1994);
   U254 : EO1 port map( A => n1946, B => n1859, C => n1898, D => n1859, Z => 
                           n2236);
   U255 : AO4 port map( A => n1983, B => n1455, C => n1878, D => n2085, Z => 
                           n2282);
   U256 : AO2 port map( A => n1914, B => n2241, C => n1916, D => n2003, Z => 
                           n2230);
   U257 : IVDA port map( A => n1902, Y => n1888, Z => n2322);
   U258 : AO2 port map( A => n1977, B => n1900, C => n2322, D => n1859, Z => 
                           n2201);
   U260 : IVDA port map( A => n1923, Y => n1455, Z => n2312);
   U261 : IVI port map( A => n2197, Z => n6747);
   U263 : AO4 port map( A => n1878, B => n1928, C => n6774, D => n1930, Z => 
                           n1925);
   U265 : AO3 port map( A => n1940, B => n1631, C => n1942, D => n1943, Z => 
                           n1939);
   U268 : AO2 port map( A => n1944, B => n2312, C => n2318, D => n1874, Z => 
                           n1943);
   U270 : EO1 port map( A => n1946, B => n1890, C => n1948, D => n6775, Z => 
                           n1942);
   U272 : IVI port map( A => n1975, Z => n6733);
   U273 : IVI port map( A => n2111, Z => n6764);
   U274 : AO6 port map( A => n6751, B => n2093, C => n2043, Z => n2085);
   U276 : IVDA port map( A => n1900, Y => n1792, Z => n2315);
   U277 : AO3 port map( A => n1998, B => n2010, C => n1890, D => n6733, Z => 
                           n2008);
   U278 : AO2 port map( A => n2000, B => n2317, C => n2319, D => n1948, Z => 
                           n2009);
   U280 : AO3 port map( A => n2083, B => n2084, C => n2313, D => n2085, Z => 
                           n2079);
   U281 : AO2 port map( A => n2317, B => n2239, C => n6738, D => n2312, Z => 
                           n2234);
   U283 : AO4 port map( A => n1888, B => n2140, C => n2048, D => n1631, Z => 
                           n2262);
   U284 : AO2 port map( A => n1914, B => n1915, C => n1916, D => n1859, Z => 
                           n1913);
   U285 : AO7 port map( A => n1978, B => n1979, C => n1980, Z => n1957);
   U286 : AO4 port map( A => n1675, B => n1983, C => n6776, D => n1972, Z => 
                           n1978);
   U288 : AO4 port map( A => n1915, B => n1878, C => n6774, D => n6750, Z => 
                           n1979);
   U290 : AO4 port map( A => n1792, B => n1874, C => n1843, D => n6730, Z => 
                           n2059);
   U291 : AO6 port map( A => n1901, B => n2126, C => n6670, Z => n2125);
   U293 : AO2 port map( A => n2115, B => n1916, C => n2129, D => n1914, Z => 
                           n2128);
   U294 : AO4 port map( A => n2055, B => n1455, C => n1843, D => n1863, Z => 
                           n2065);
   U295 : AO2 port map( A => n2054, B => n2322, C => n2055, D => n2312, Z => 
                           n2053);
   U296 : AO2 port map( A => n2318, B => n1944, C => n2319, D => n2118, Z => 
                           n2180);
   U297 : EON1 port map( A => n1878, B => n2102, C => n2241, D => n2318, Z => 
                           n2261);
   U298 : AO6 port map( A => n6769, B => n6765, C => n1455, Z => n1855);
   U299 : AO2 port map( A => n2318, B => n1930, C => n2319, D => n2129, Z => 
                           n2202);
   U300 : ND4 port map( A => n1992, B => n1993, C => n1994, D => n1995, Z => 
                           n1991);
   U301 : AO2 port map( A => n2000, B => n2312, C => n2319, D => n6745, Z => 
                           n1993);
   U302 : EO1 port map( A => n2002, B => n2315, C => n2003, D => n1888, Z => 
                           n1992);
   U303 : ND4 port map( A => n6742, B => n2275, C => n2276, D => n2277, Z => 
                           n2266);
   U304 : AO2 port map( A => n2315, B => n6747, C => n6732, D => n2317, Z => 
                           n2275);
   U305 : AO2 port map( A => n2048, B => n2318, C => n2319, D => n6751, Z => 
                           n2276);
   U306 : AO6 port map( A => n2313, B => n1890, C => n2151, Z => n2199);
   U307 : AO2 port map( A => n2178, B => n2315, C => n2322, D => n2032, Z => 
                           n2171);
   U308 : AO7 port map( A => n1940, B => n2188, C => n2313, Z => n2185);
   U309 : AO7 port map( A => n6748, B => n6776, C => n2184, Z => n2166);
   U310 : IVDA port map( A => n166, Y => n1876, Z => n2304);
   U311 : AO6 port map( A => n2029, B => n2030, C => n4558, Z => n2015);
   U312 : AO2 port map( A => n1914, B => n1928, C => n6737, D => n1916, Z => 
                           n2030);
   U313 : AO2 port map( A => n1901, B => n2033, C => n2034, D => n2320, Z => 
                           n2029);
   U314 : AO7 port map( A => n2052, B => n2311, C => n2053, Z => n2033);
   U315 : ND4 port map( A => n2035, B => n2036, C => n2037, D => n2038, Z => 
                           n2034);
   U316 : AO2 port map( A => n2042, B => n2311, C => n2043, D => n2313, Z => 
                           n2037);
   U317 : AO2 port map( A => n2319, B => n2049, C => n1935, D => n2315, Z => 
                           n2035);
   U318 : IVI port map( A => n1937, Z => n6774);
   U319 : IVI port map( A => n1924, Z => n6776);
   U320 : NR4 port map( A => n2086, B => n2087, C => n2088, D => n2089, Z => 
                           n2070);
   U321 : AO4 port map( A => n1843, B => n1936, C => n2316, D => n1888, Z => 
                           n2088);
   U322 : AO4 port map( A => n1859, B => n6776, C => n1455, D => n2090, Z => 
                           n2089);
   U323 : AO4 port map( A => n6731, B => n6775, C => n6774, D => n2092, Z => 
                           n2086);
   U324 : IVDA port map( A => n1881, Y => n1631, Z => n2319);
   U325 : AO3 port map( A => n6776, B => n2078, C => n2079, D => n2080, Z => 
                           n2074);
   U326 : AO4 port map( A => n6731, B => n1843, C => n1631, D => n2077, Z => 
                           n2075);
   U327 : IVDA port map( A => n2044, Y => n1878, Z => n2313);
   U328 : AO2 port map( A => n2081, B => n2082, C => n1998, D => n6764, Z => 
                           n2080);
   U329 : AO4 port map( A => n6755, B => n1888, C => n6768, D => n1847, Z => 
                           n2082);
   U330 : AO3 port map( A => n6776, B => n6761, C => n2256, D => n2257, Z => 
                           n2254);
   U331 : ND3 port map( A => n6733, B => n2313, C => n1859, Z => n2256);
   U332 : EO1 port map( A => n2310, B => n2115, C => n6774, D => n1915, Z => 
                           n2257);
   U334 : AO7 port map( A => n1919, B => n2311, C => n1920, Z => n1918);
   U335 : AO2 port map( A => n6737, B => n2322, C => n6735, D => n2312, Z => 
                           n1920);
   U336 : AO7 port map( A => n1901, B => n2251, C => n2252, Z => n2250);
   U337 : NR4 port map( A => n2260, B => n2261, C => n2262, D => n2263, Z => 
                           n2251);
   U338 : AO2 port map( A => n1980, B => n2253, C => n2184, D => n2254, Z => 
                           n2252);
   U339 : AO4 port map( A => n2316, B => n1455, C => n2002, D => n1843, Z => 
                           n2263);
   U340 : ND4 port map( A => n1960, B => n1961, C => n6736, D => n1963, Z => 
                           n1959);
   U341 : AO2 port map( A => n2321, B => n1900, C => n1977, D => n2317, Z => 
                           n1960);
   U342 : AO2 port map( A => n2318, B => n6758, C => n1975, D => n2319, Z => 
                           n1961);
   U343 : IVDA port map( A => n1945, Y => n1847, Z => n2318);
   U344 : AO4 port map( A => n1888, B => n1948, C => n2316, D => n1792, Z => 
                           n2005);
   U345 : AO3 port map( A => n2007, B => n1847, C => n2008, D => n2009, Z => 
                           n2004);
   U346 : AO4 port map( A => n1843, B => n2114, C => n1888, D => n2115, Z => 
                           n2113);
   U347 : AO2 port map( A => n2318, B => n2118, C => n4562, D => n1900, Z => 
                           n2116);
   U348 : IVDA port map( A => n1934, Y => n1843, Z => n2317);
   U349 : AO2 port map( A => n1938, B => n2317, C => n2318, D => n2140, Z => 
                           n2139);
   U350 : AO7 port map( A => n1894, B => n1675, C => n2258, Z => n2253);
   U352 : AO2 port map( A => n6738, B => n2259, C => n1924, D => n2077, Z => 
                           n2258);
   U353 : AO7 port map( A => n1587, B => n1909, C => n6774, Z => n2259);
   U354 : AO3 port map( A => n6773, B => n1869, C => n1870, D => n1871, Z => 
                           n1854);
   U355 : AO4 port map( A => n2000, B => n1631, C => n2314, D => n1898, Z => 
                           n2019);
   U356 : AO3 port map( A => n6775, B => n2049, C => n2226, D => n2227, Z => 
                           n2212);
   U357 : AO2 port map( A => n2000, B => n2105, C => n2319, D => n6760, Z => 
                           n2227);
   U358 : EO1 port map( A => n2228, B => n1924, C => n2155, D => n6773, Z => 
                           n2226);
   U359 : NR3 port map( A => n2135, B => n2136, C => n2137, Z => n2124);
   U360 : AO4 port map( A => n1455, B => n6745, C => n2316, D => n1888, Z => 
                           n2137);
   U361 : AO3 port map( A => n6775, B => n1889, C => n2138, D => n2139, Z => 
                           n2135);
   U362 : AO4 port map( A => n2055, B => n1792, C => n2054, D => n1631, Z => 
                           n2136);
   U363 : AO6 port map( A => n2232, B => n2320, C => n2508, Z => n2231);
   U364 : ND4 port map( A => n2234, B => n2235, C => n2236, D => n2237, Z => 
                           n2232);
   U365 : AO2 port map( A => n2141, B => n6777, C => n2315, D => n2238, Z => 
                           n2237);
   U366 : AO6 port map( A => n2142, B => n2320, C => n2143, Z => n2120);
   U367 : AO4 port map( A => n2144, B => n6779, C => n2145, D => n6780, Z => 
                           n2143);
   U368 : AO3 port map( A => n1843, B => n2155, C => n2156, D => n2157, Z => 
                           n2142);
   U369 : NR4 port map( A => n1763, B => n1587, C => n2321, D => n6770, Z => 
                           n2207);
   U370 : AO4 port map( A => n1455, B => n6769, C => n2208, D => n1843, Z => 
                           n2206);
   U371 : AO3 port map( A => n6776, B => n6750, C => n2132, D => n2133, Z => 
                           n2131);
   U373 : AO2 port map( A => n2083, B => n2313, C => n2084, D => n2310, Z => 
                           n2132);
   U374 : AO6 port map( A => n1937, B => n1973, C => n1873, Z => n2133);
   U375 : AO7 port map( A => n1901, B => n2190, C => n2191, Z => n2189);
   U377 : AO2 port map( A => n1980, B => n2192, C => n2184, D => n2193, Z => 
                           n2191);
   U378 : AO3 port map( A => n1587, B => n6749, C => n2199, D => n2200, Z => 
                           n2192);
   U379 : AO6 port map( A => n1858, B => n2321, C => n2208, Z => n2002);
   U380 : NR3 port map( A => n1859, B => n1587, C => n6772, Z => n2010);
   U381 : AO4 port map( A => n1878, B => n6671, C => n1940, D => n6776, Z => 
                           n1987);
   U382 : AO4 port map( A => n1878, B => n6764, C => n1675, D => n6733, Z => 
                           n2148);
   U383 : AO7 port map( A => n6774, B => n1874, C => n6672, Z => n2149);
   U384 : AO4 port map( A => n1792, B => n6754, C => n1888, D => n6760, Z => 
                           n2225);
   U385 : AO2 port map( A => n1924, B => n1930, C => n6732, D => n2313, Z => 
                           n2219);
   U386 : AO6 port map( A => n6754, B => n1864, C => n1843, Z => n2273);
   U387 : AO2 port map( A => n2141, B => n1937, C => n1946, D => n2314, Z => 
                           n2138);
   U388 : AO3 port map( A => n6731, B => n2194, C => n2195, D => n2196, Z => 
                           n2193);
   U389 : AO7 port map( A => n1975, B => n2197, C => n2313, Z => n2195);
   U390 : AO6 port map( A => n2198, B => n1587, C => n1924, Z => n2194);
   U391 : AO4 port map( A => n1857, B => n1888, C => n1843, D => n1860, Z => 
                           n1856);
   U392 : AO3 port map( A => n2305, B => n1843, C => n2026, D => n2027, Z => 
                           n2017);
   U393 : AO2 port map( A => n2318, B => n6733, C => n1900, D => n6734, Z => 
                           n2027);
   U394 : AO4 port map( A => n2061, B => n1936, C => n2062, D => n1888, Z => 
                           n2060);
   U395 : AO6 port map( A => n2310, B => n2049, C => n2152, Z => n2144);
   U396 : AO4 port map( A => n1887, B => n6776, C => n6731, D => n2153, Z => 
                           n2152);
   U397 : AO6 port map( A => n2154, B => n2321, C => n1937, Z => n2153);
   U398 : AO2 port map( A => n1763, B => n2215, C => n2216, D => n1873, Z => 
                           n2214);
   U399 : AO3 port map( A => n1878, B => n1970, C => n2222, D => n2223, Z => 
                           n2215);
   U400 : AO3 port map( A => n6774, B => n6744, C => n2218, D => n2219, Z => 
                           n2216);
   U401 : AO2 port map( A => n1901, B => n2168, C => n2169, D => n2320, Z => 
                           n2167);
   U402 : AO3 port map( A => n2054, B => n1843, C => n2179, D => n2180, Z => 
                           n2168);
   U403 : ND3 port map( A => n2170, B => n2171, C => n2172, Z => n2169);
   U404 : AO3 port map( A => n6731, B => n1455, C => n2270, D => n2271, Z => 
                           n2269);
   U405 : AO2 port map( A => n1900, B => n2090, C => n2111, D => n2322, Z => 
                           n2270);
   U406 : AO6 port map( A => n2305, B => n6755, C => n2051, Z => n1935);
   U407 : AO2 port map( A => n1924, B => n1889, C => n2028, D => n2310, Z => 
                           n2200);
   U408 : AO2 port map( A => n2310, B => n6758, C => n1937, D => n2119, Z => 
                           n2223);
   U409 : AO2 port map( A => n2321, B => n2317, C => n2312, D => n1936, Z => 
                           n2170);
   U410 : AO2 port map( A => n2322, B => n6751, C => n2316, D => n2312, Z => 
                           n2130);
   U411 : AO6 port map( A => n2305, B => n1763, C => n2024, Z => n2081);
   U412 : AO7 port map( A => n2011, B => n2187, C => n2310, Z => n2186);
   U413 : AO7 port map( A => n226, B => n2391, C => n6790, Z => n171);
   U414 : NR3 port map( A => n1876, B => n156, C => n157, Z => n226);
   U415 : AO7 port map( A => n66, B => n153, C => n67, Z => n149);
   U416 : AO7 port map( A => n66, B => n112, C => n67, Z => n108);
   U417 : AO7 port map( A => n66, B => n62, C => n67, Z => n57);
   U418 : IVDA port map( A => n63, Y => n1904, Z => n2325);
   U419 : OR3 port map( A => n153, B => n2325, C => n6782, Z => n121);
   U421 : OR3 port map( A => n112, B => n2325, C => n6784, Z => n80);
   U422 : OR3 port map( A => n62, B => n2325, C => n2504, Z => n21);
   U423 : AO4 port map( A => n1877, B => n68, C => n6795, D => n252, Z => n157)
                           ;
   U424 : IVDA port map( A => n324, Y => n2066, Z => n2326);
   U425 : NR3 port map( A => v_CALCULATION_CNTR_1_port, B => n2255, C => n6793,
                           Z => n225);
   U426 : AO4 port map( A => CE_I, B => n2181, C => n1848, D => n2391, Z => 
                           n4596);
   U427 : NR4 port map( A => n1853, B => n1854, C => n1855, D => n1856, Z => 
                           n1852);
   U428 : AO3 port map( A => n1901, B => n1911, C => n1912, D => n1913, Z => 
                           n1849);
   U429 : AO4 port map( A => CE_I, B => n2217, C => n2012, D => n2391, Z => 
                           n4598);
   U430 : NR3 port map( A => n2017, B => n2018, C => n2019, Z => n2016);
   U431 : IVDA port map( A => n1927, Y => n1675, Z => n2310);
   U432 : IVDA port map( A => n2020, Y => n1903, Z => n2314);
   U433 : EO1 port map( A => n2039, B => n2040, C => n1985, D => n1873, Z => 
                           n2038);
   U434 : AO4 port map( A => n1969, B => n1455, C => n6768, D => n1888, Z => 
                           n2040);
   U435 : AO2 port map( A => n2096, B => n2308, C => n1587, D => n2097, Z => 
                           n2095);
   U436 : AO3 port map( A => n6778, B => n2106, C => n2107, D => n2108, Z => 
                           n2096);
   U437 : AO3 port map( A => n6778, B => n1903, C => n1870, D => n2099, Z => 
                           n2097);
   U438 : NR4 port map( A => n1891, B => n1892, C => n1850, D => n2320, Z => 
                           n1851);
   U439 : AO4 port map( A => n1894, B => n1455, C => n1895, D => n1843, Z => 
                           n1892);
   U440 : AO3 port map( A => n1896, B => n1897, C => n1898, D => n1899, Z => 
                           n1891);
   U441 : AO2 port map( A => n2315, B => n1889, C => n2322, D => n6754, Z => 
                           n1899);
   U442 : AO4 port map( A => CE_I, B => n2220, C => n2067, D => n2391, Z => 
                           n4599);
   U443 : AO6 port map( A => n1901, B => n2068, C => n2069, Z => n2067);
   U444 : AO4 port map( A => n2070, B => n4560, C => n2071, D => n2072, Z => 
                           n2069);
   U445 : AO4 port map( A => n2094, B => n1850, C => n4558, D => n2095, Z => 
                           n2068);
   U446 : AO2 port map( A => n2100, B => n1897, C => n6767, D => n6777, Z => 
                           n2099);
   U447 : AO3 port map( A => n6755, B => n6771, C => n6756, D => n2104, Z => 
                           n2100);
   U448 : AO4 port map( A => n1878, B => n2058, C => n6774, D => n2032, Z => 
                           n2056);
   U449 : AO6 port map( A => n6671, B => n1970, C => n2308, Z => n2057);
   U450 : AO7 port map( A => CE_I, B => n2205, C => n1950, Z => n4597);
   U451 : AO2 port map( A => n1951, B => n1952, C => n1953, D => n1954, Z => 
                           n1950);
   U452 : AO7 port map( A => n1990, B => n2320, C => n1991, Z => n1952);
   U453 : AO3 port map( A => n1955, B => n6779, C => n1957, D => n1958, Z => 
                           n1954);
   U454 : AO3 port map( A => CE_I, B => n2240, C => n2248, D => n2249, Z => 
                           n4603);
   U455 : ND4 port map( A => n1953, B => n2266, C => n2267, D => n2268, Z => 
                           n2248);
   U456 : AO2 port map( A => n6741, B => n1914, C => n2246, D => n1916, Z => 
                           n2267);
   U457 : AO2 port map( A => n1885, B => n2317, C => n2322, D => n1935, Z => 
                           n1933);
   U458 : AO2 port map( A => n1936, B => n2315, C => n1937, D => n1938, Z => 
                           n1932);
   U459 : AO4 port map( A => n266, B => n6789, C => n6793, D => n2298, Z => 
                           n153);
   U460 : AO4 port map( A => n6786, B => n6793, C => n2255, D => n2300, Z => 
                           n112);
   U461 : AO7 port map( A => n1885, B => n1455, C => n2247, Z => n2242);
   U462 : AO4 port map( A => n1888, B => n6739, C => n2308, D => n2245, Z => 
                           n2243);
   U463 : EO1 port map( A => n2314, B => n1900, C => n2090, D => n1843, Z => 
                           n2247);
   U465 : IVDA port map( A => n2006, Y => n1889, Z => n2316);
   U466 : IVDA port map( A => n1976, Y => n1890, Z => n2321);
   U467 : AO3 port map( A => n1878, B => n6733, C => n2045, D => n2046, Z => 
                           n2042);
   U468 : AO2 port map( A => n2322, B => n1964, C => n2312, D => n1965, Z => 
                           n1963);
   U469 : AO7 port map( A => n1858, B => n1969, C => n1970, Z => n1964);
   U470 : NR4 port map( A => n1850, B => n2064, C => n2320, D => n2065, Z => 
                           n2013);
   U471 : AO4 port map( A => n1631, B => n6764, C => n4562, D => n1847, Z => 
                           n2064);
   U472 : EO1 port map( A => n1946, B => n1969, C => n6775, D => n2054, Z => 
                           n2117);
   U473 : AO3 port map( A => CE_I, B => n2233, C => n2163, D => n2164, Z => 
                           n4601);
   U474 : AO3 port map( A => n2165, B => n2166, C => n1951, D => n2167, Z => 
                           n2164);
   U475 : AO3 port map( A => n1887, B => n6752, C => n2185, D => n2186, Z => 
                           n2165);
   U476 : AO3 port map( A => CE_I, B => n2183, C => n2209, D => n2210, Z => 
                           n4602);
   U477 : AO3 port map( A => n2229, B => n1893, C => n2230, D => n2231, Z => 
                           n2209);
   U478 : AO4 port map( A => n2212, B => n2213, C => n1901, D => n2214, Z => 
                           n2211);
   U479 : AO3 port map( A => n1969, B => n1898, C => n2264, D => n2265, Z => 
                           n2260);
   U480 : AO7 port map( A => n2187, B => n2051, C => n2315, Z => n2265);
   U481 : ND4 port map( A => v_CALCULATION_CNTR_1_port, B => n2301, C => n2255,
                           D => n1877, Z => n2303);
   U482 : AO4 port map( A => n1847, B => n2073, C => n6774, D => n2102, Z => 
                           n2173);
   U483 : AO4 port map( A => n6771, B => n6752, C => n1985, D => n2176, Z => 
                           n2174);
   U484 : IVDA port map( A => n1873, Y => n1763, Z => n2311);
   U485 : AO2 port map( A => n2318, B => n6735, C => n2319, D => n1969, Z => 
                           n2235);
   U486 : AO3 port map( A => n1792, B => n6730, C => n1879, D => n1880, Z => 
                           n1853);
   U487 : AO6 port map( A => n2319, B => n6751, C => n4560, Z => n1880);
   U488 : AO2 port map( A => n1884, B => n1885, C => n1886, D => n1887, Z => 
                           n1879);
   U489 : AO7 port map( A => n1878, B => n6772, C => n1847, Z => n1884);
   U490 : AO3 port map( A => n2021, B => n1897, C => n2022, D => n6753, Z => 
                           n2018);
   U491 : AO6 port map( A => n1890, B => n2311, C => n2024, Z => n2021);
   U492 : ND3 port map( A => n6764, B => n1859, C => n2312, Z => n2022);
   U493 : IVDA port map( A => n2025, Y => n1858, Z => n2305);
   U494 : AO2 port map( A => n2109, B => n1897, C => n6768, D => n2093, Z => 
                           n2108);
   U495 : AO3 port map( A => n1763, B => n6747, C => n2110, D => n6771, Z => 
                           n2109);
   U496 : AO7 port map( A => n2111, B => n2316, C => n1763, Z => n2110);
   U497 : AO3 port map( A => n2308, B => n2160, C => n1873, D => n6743, Z => 
                           n2156);
   U498 : AO4 port map( A => n2106, B => n6774, C => n2077, D => n1878, Z => 
                           n2162);
   U499 : IVDA port map( A => n1893, Y => n1901, Z => n2320);
   U500 : AO7 port map( A => v_CALCULATION_CNTR_2_port, B => n230, C => n1904, 
                           Z => n156);
   U501 : NR4 port map( A => n2255, B => n6795, C => n1877, D => 
                           v_CALCULATION_CNTR_1_port, Z => n290);
   U502 : AO4 port map( A => v_CALCULATION_CNTR_2_port, B => n68, C => n1882, D
                           => n70, Z => n62);
   U503 : EO1 port map( A => n2497, B => n2498, C => n68, D => n1877, Z => 
                           n2496);
   U504 : AO7 port map( A => n262, B => n2391, C => n240, Z => n254);
   U505 : AO6 port map( A => n264, B => n1877, C => n2325, Z => n262);
   U506 : AO7 port map( A => n267, B => n230, C => n6795, Z => n264);
   U507 : AO7 port map( A => n290, B => n155, C => n67, Z => n287);
   U509 : AO4 port map( A => CE_I, B => n1947, C => n336, D => n2391, Z => 
                           n4564);
   U510 : ND4 port map( A => n391, B => n392, C => n393, D => n394, Z => n337);
   U511 : ND4 port map( A => n339, B => n340, C => n341, D => n342, Z => n338);
   U512 : AO4 port map( A => CE_I, B => n1929, C => n444, D => n2391, Z => 
                           n4565);
   U513 : ND4 port map( A => n467, B => n468, C => n469, D => n470, Z => n445);
   U514 : ND4 port map( A => n447, B => n448, C => n449, D => n450, Z => n446);
   U515 : AO4 port map( A => CE_I, B => n1867, C => n488, D => n2391, Z => 
                           n4566);
   U516 : ND4 port map( A => n511, B => n512, C => n513, D => n514, Z => n489);
   U517 : ND4 port map( A => n491, B => n492, C => n493, D => n494, Z => n490);
   U518 : AO4 port map( A => CE_I, B => n1981, C => n532, D => n2391, Z => 
                           n4567);
   U519 : ND4 port map( A => n555, B => n556, C => n557, D => n558, Z => n533);
   U520 : ND4 port map( A => n535, B => n536, C => n537, D => n538, Z => n534);
   U521 : AO4 port map( A => CE_I, B => n1974, C => n576, D => n2391, Z => 
                           n4568);
   U522 : ND4 port map( A => n599, B => n600, C => n601, D => n602, Z => n577);
   U523 : ND4 port map( A => n579, B => n580, C => n581, D => n582, Z => n578);
   U524 : AO4 port map( A => CE_I, B => n1949, C => n620, D => n2391, Z => 
                           n4569);
   U525 : ND4 port map( A => n643, B => n644, C => n645, D => n646, Z => n621);
   U526 : ND4 port map( A => n623, B => n624, C => n625, D => n626, Z => n622);
   U527 : AO4 port map( A => CE_I, B => n1989, C => n664, D => n2391, Z => 
                           n4570);
   U528 : ND4 port map( A => n687, B => n688, C => n689, D => n690, Z => n665);
   U529 : ND4 port map( A => n667, B => n668, C => n669, D => n670, Z => n666);
   U530 : AO4 port map( A => CE_I, B => n1966, C => n708, D => n2391, Z => 
                           n4571);
   U531 : ND4 port map( A => n731, B => n732, C => n733, D => n734, Z => n709);
   U532 : ND4 port map( A => n711, B => n712, C => n713, D => n714, Z => n710);
   U533 : AO4 port map( A => CE_I, B => n1922, C => n752, D => n2391, Z => 
                           n4572);
   U534 : ND4 port map( A => n775, B => n776, C => n777, D => n778, Z => n753);
   U535 : ND4 port map( A => n755, B => n756, C => n757, D => n758, Z => n754);
   U536 : AO4 port map( A => CE_I, B => n1956, C => n796, D => n2391, Z => 
                           n4573);
   U537 : ND4 port map( A => n819, B => n820, C => n821, D => n822, Z => n797);
   U538 : ND4 port map( A => n799, B => n800, C => n801, D => n802, Z => n798);
   U539 : AO4 port map( A => CE_I, B => n1999, C => n840, D => n2391, Z => 
                           n4574);
   U540 : ND4 port map( A => n863, B => n864, C => n865, D => n866, Z => n841);
   U541 : ND4 port map( A => n843, B => n844, C => n845, D => n846, Z => n842);
   U542 : AO4 port map( A => CE_I, B => n1968, C => n884, D => n2391, Z => 
                           n4575);
   U543 : ND4 port map( A => n907, B => n908, C => n909, D => n910, Z => n885);
   U544 : ND4 port map( A => n887, B => n888, C => n889, D => n890, Z => n886);
   U545 : AO4 port map( A => CE_I, B => n1872, C => n928, D => n2391, Z => 
                           n4576);
   U546 : ND4 port map( A => n951, B => n952, C => n953, D => n954, Z => n929);
   U547 : ND4 port map( A => n931, B => n932, C => n933, D => n934, Z => n930);
   U548 : AO4 port map( A => CE_I, B => n1962, C => n972, D => n2391, Z => 
                           n4577);
   U549 : ND4 port map( A => n995, B => n996, C => n997, D => n998, Z => n973);
   U550 : ND4 port map( A => n975, B => n976, C => n977, D => n978, Z => n974);
   U551 : AO4 port map( A => CE_I, B => n1868, C => n1016, D => n2391, Z => 
                           n4578);
   U553 : ND4 port map( A => n1039, B => n1040, C => n1041, D => n1042, Z => 
                           n1017);
   U554 : ND4 port map( A => n1019, B => n1020, C => n1021, D => n1022, Z => 
                           n1018);
   U555 : AO4 port map( A => CE_I, B => n2001, C => n1060, D => n2391, Z => 
                           n4579);
   U556 : ND4 port map( A => n1083, B => n1084, C => n1085, D => n1086, Z => 
                           n1061);
   U557 : ND4 port map( A => n1063, B => n1064, C => n1065, D => n1066, Z => 
                           n1062);
   U558 : AO4 port map( A => CE_I, B => n1982, C => n1104, D => n2391, Z => 
                           n4580);
   U559 : ND4 port map( A => n1127, B => n1128, C => n1129, D => n1130, Z => 
                           n1105);
   U560 : ND4 port map( A => n1107, B => n1108, C => n1109, D => n1110, Z => 
                           n1106);
   U561 : AO4 port map( A => CE_I, B => n1984, C => n1148, D => n2391, Z => 
                           n4581);
   U562 : ND4 port map( A => n1171, B => n1172, C => n1173, D => n1174, Z => 
                           n1149);
   U563 : ND4 port map( A => n1151, B => n1152, C => n1153, D => n1154, Z => 
                           n1150);
   U564 : AO4 port map( A => CE_I, B => n1967, C => n1192, D => n2391, Z => 
                           n4582);
   U565 : ND4 port map( A => n1215, B => n1216, C => n1217, D => n1218, Z => 
                           n1193);
   U566 : ND4 port map( A => n1195, B => n1196, C => n1197, D => n1198, Z => 
                           n1194);
   U567 : AO4 port map( A => CE_I, B => n2023, C => n1236, D => n2391, Z => 
                           n4583);
   U568 : ND4 port map( A => n1259, B => n1260, C => n1261, D => n1262, Z => 
                           n1237);
   U569 : ND4 port map( A => n1239, B => n1240, C => n1241, D => n1242, Z => 
                           n1238);
   U570 : AO4 port map( A => CE_I, B => n1905, C => n1280, D => n2391, Z => 
                           n4584);
   U571 : ND4 port map( A => n1303, B => n1304, C => n1305, D => n1306, Z => 
                           n1281);
   U572 : ND4 port map( A => n1283, B => n1284, C => n1285, D => n1286, Z => 
                           n1282);
   U573 : AO4 port map( A => CE_I, B => n1931, C => n1324, D => n2391, Z => 
                           n4585);
   U574 : ND4 port map( A => n1347, B => n1348, C => n1349, D => n1350, Z => 
                           n1325);
   U575 : ND4 port map( A => n1327, B => n1328, C => n1329, D => n1330, Z => 
                           n1326);
   U576 : AO4 port map( A => CE_I, B => n1921, C => n1368, D => n2391, Z => 
                           n4586);
   U577 : ND4 port map( A => n1391, B => n1392, C => n1393, D => n1394, Z => 
                           n1369);
   U578 : ND4 port map( A => n1371, B => n1372, C => n1373, D => n1374, Z => 
                           n1370);
   U579 : AO4 port map( A => CE_I, B => n1906, C => n1412, D => n2391, Z => 
                           n4587);
   U580 : ND4 port map( A => n1435, B => n1436, C => n1437, D => n1438, Z => 
                           n1413);
   U581 : ND4 port map( A => n1415, B => n1416, C => n1417, D => n1418, Z => 
                           n1414);
   U582 : AO4 port map( A => CE_I, B => n1862, C => n1456, D => n2391, Z => 
                           n4588);
   U583 : ND4 port map( A => n1479, B => n1480, C => n1481, D => n1482, Z => 
                           n1457);
   U584 : ND4 port map( A => n1459, B => n1460, C => n1461, D => n1462, Z => 
                           n1458);
   U585 : AO4 port map( A => CE_I, B => n1910, C => n1500, D => n2391, Z => 
                           n4589);
   U586 : ND4 port map( A => n1523, B => n1524, C => n1525, D => n1526, Z => 
                           n1501);
   U587 : ND4 port map( A => n1503, B => n1504, C => n1505, D => n1506, Z => 
                           n1502);
   U588 : AO4 port map( A => CE_I, B => n1865, C => n1544, D => n2391, Z => 
                           n4590);
   U589 : ND4 port map( A => n1567, B => n1568, C => n1569, D => n1570, Z => 
                           n1545);
   U590 : ND4 port map( A => n1547, B => n1548, C => n1549, D => n1550, Z => 
                           n1546);
   U591 : AO4 port map( A => CE_I, B => n1861, C => n1588, D => n2391, Z => 
                           n4591);
   U592 : ND4 port map( A => n1611, B => n1612, C => n1613, D => n1614, Z => 
                           n1589);
   U593 : ND4 port map( A => n1591, B => n1592, C => n1593, D => n1594, Z => 
                           n1590);
   U594 : AO4 port map( A => CE_I, B => n1908, C => n1632, D => n2391, Z => 
                           n4592);
   U595 : ND4 port map( A => n1655, B => n1656, C => n1657, D => n1658, Z => 
                           n1633);
   U597 : ND4 port map( A => n1635, B => n1636, C => n1637, D => n1638, Z => 
                           n1634);
   U598 : AO4 port map( A => CE_I, B => n1917, C => n1676, D => n2391, Z => 
                           n4593);
   U599 : ND4 port map( A => n1699, B => n1700, C => n1701, D => n1702, Z => 
                           n1677);
   U600 : ND4 port map( A => n1679, B => n1680, C => n1681, D => n1682, Z => 
                           n1678);
   U601 : AO4 port map( A => CE_I, B => n1941, C => n1720, D => n2391, Z => 
                           n4594);
   U602 : ND4 port map( A => n1743, B => n1744, C => n1745, D => n1746, Z => 
                           n1721);
   U603 : ND4 port map( A => n1723, B => n1724, C => n1725, D => n1726, Z => 
                           n1722);
   U604 : AO4 port map( A => CE_I, B => n1866, C => n1764, D => n2391, Z => 
                           n4595);
   U605 : ND4 port map( A => n1809, B => n1810, C => n1811, D => n1812, Z => 
                           n1765);
   U606 : ND4 port map( A => n1767, B => n1768, C => n1769, D => n1770, Z => 
                           n1766);
   U607 : EON1 port map( A => n1833, B => n6788, C => n1833, D => n287, Z => 
                           n6728);
   U608 : NR4 port map( A => n2031, B => n65, C => n290, D => n6805, Z => n2499
                           );
   U609 : NR3 port map( A => i_SRAM_ADDR_WR02, B => n2480, C => 
                           i_SRAM_ADDR_WR01, Z => n2471);
   U610 : IVDA port map( A => n292, Y => n2041, Z => n2324);
   U611 : NR3 port map( A => n6803, B => n1832, C => n1719, Z => n292);
   U612 : AN3 port map( A => n1832, B => n1719, C => n312, Z => n324);
   U613 : AO4 port map( A => n268, B => n2031, C => n2479, D => n271, Z => 
                           n6723);
   U614 : IVDA port map( A => n304, Y => n2076, Z => n2323);
   U615 : ND2I port map( A => n2293, B => n2294, Z => n1969);
   U616 : AO2 port map( A => v_TEMP_VECTOR_28_port, B => n112, C => 
                           v_TEMP_VECTOR_20_port, D => n153, Z => n2294);
   U617 : AO2 port map( A => v_TEMP_VECTOR_12_port, B => n1876, C => 
                           v_TEMP_VECTOR_4_port, D => n2281, Z => n2293);
   U618 : ND2I port map( A => n2285, B => n2286, Z => n1897);
   U619 : AO2 port map( A => v_TEMP_VECTOR_31_port, B => n112, C => 
                           v_TEMP_VECTOR_23_port, D => n153, Z => n2286);
   U620 : AO2 port map( A => v_TEMP_VECTOR_15_port, B => n1876, C => 
                           v_TEMP_VECTOR_7_port, D => n2281, Z => n2285);
   U621 : NR3 port map( A => v_CALCULATION_CNTR_7_port, B => 
                           v_CALCULATION_CNTR_6_port, C => 
                           v_CALCULATION_CNTR_5_port, Z => n2306);
   U622 : ND3 port map( A => n2306, B => n1844, C => v_CALCULATION_CNTR_3_port,
                           Z => n230);
   U623 : AO2 port map( A => v_TEMP_VECTOR_27_port, B => n112, C => 
                           v_TEMP_VECTOR_19_port, D => n153, Z => n2292);
   U624 : AO2 port map( A => v_TEMP_VECTOR_11_port, B => n1876, C => 
                           v_TEMP_VECTOR_3_port, D => n2281, Z => n2291);
   U625 : IVDA port map( A => n2047, Y => n1587, Z => n2308);
   U626 : AO2 port map( A => v_TEMP_VECTOR_29_port, B => n112, C => 
                           v_TEMP_VECTOR_21_port, D => n153, Z => n2288);
   U627 : AO2 port map( A => v_TEMP_VECTOR_13_port, B => n1876, C => 
                           v_TEMP_VECTOR_5_port, D => n2281, Z => n2287);
   U628 : AO3 port map( A => n2120, B => n4559, C => n2122, D => n2123, Z => 
                           n4600);
   U629 : AO3 port map( A => n1901, B => n2124, C => n1951, D => n2125, Z => 
                           n2122);
   U630 : AO2 port map( A => v_TEMP_VECTOR_26_port, B => n112, C => 
                           v_TEMP_VECTOR_18_port, D => n153, Z => n2284);
   U631 : AO2 port map( A => v_TEMP_VECTOR_10_port, B => n1876, C => 
                           v_TEMP_VECTOR_2_port, D => n2281, Z => n2283);
   U632 : AO2 port map( A => v_TEMP_VECTOR_25_port, B => n112, C => 
                           v_TEMP_VECTOR_17_port, D => n153, Z => n2290);
   U633 : AO2 port map( A => v_TEMP_VECTOR_9_port, B => n1876, C => 
                           v_TEMP_VECTOR_1_port, D => n2281, Z => n2289);
   U634 : AO2 port map( A => v_TEMP_VECTOR_30_port, B => n112, C => 
                           v_TEMP_VECTOR_22_port, D => n153, Z => n2280);
   U635 : AO2 port map( A => v_TEMP_VECTOR_14_port, B => n1876, C => 
                           v_TEMP_VECTOR_6_port, D => n2281, Z => n2279);
   U636 : AO7 port map( A => n2103, B => n171, C => n218, Z => n6709);
   U637 : AO2 port map( A => n164, B => n219, C => v_KEY32_IN_0_port, D => n162
                           , Z => n218);
   U638 : AO4 port map( A => n174, B => n220, C => n2304, D => n2181, Z => n219
                           );
   U639 : AO2 port map( A => n176, B => n221, C => n2325, D => n222, Z => n220)
                           ;
   U641 : AO3 port map( A => n159, B => n210, C => n211, D => n212, Z => n6708)
                           ;
   U642 : AO2 port map( A => v_KEY32_IN_1_port, B => n162, C => n6785, D => 
                           v_TEMP_VECTOR_1_port, Z => n212);
   U643 : AO3 port map( A => n202, B => n159, C => n203, D => n204, Z => n6707)
                           ;
   U644 : AO2 port map( A => v_KEY32_IN_2_port, B => n162, C => n6785, D => 
                           v_TEMP_VECTOR_2_port, Z => n204);
   U645 : AO3 port map( A => n159, B => n194, C => n195, D => n196, Z => n6706)
                           ;
   U646 : AO2 port map( A => v_KEY32_IN_3_port, B => n162, C => n6785, D => 
                           v_TEMP_VECTOR_3_port, Z => n196);
   U647 : AO3 port map( A => n159, B => n188, C => n189, D => n190, Z => n6705)
                           ;
   U648 : AO2 port map( A => v_KEY32_IN_4_port, B => n162, C => n6785, D => 
                           v_TEMP_VECTOR_4_port, Z => n190);
   U649 : AO3 port map( A => n181, B => n159, C => n182, D => n183, Z => n6704)
                           ;
   U650 : AO2 port map( A => v_KEY32_IN_5_port, B => n162, C => n6785, D => 
                           v_TEMP_VECTOR_5_port, Z => n183);
   U651 : AO7 port map( A => n2121, B => n171, C => n172, Z => n6703);
   U652 : AO2 port map( A => n164, B => n173, C => v_KEY32_IN_6_port, D => n162
                           , Z => n172);
   U653 : AO4 port map( A => n2304, B => n2183, C => n174, D => n175, Z => n173
                           );
   U654 : AO2 port map( A => n176, B => n177, C => n2325, D => n178, Z => n175)
                           ;
   U655 : AO3 port map( A => n158, B => n159, C => n160, D => n161, Z => n6702)
                           ;
   U656 : AO2 port map( A => v_KEY32_IN_7_port, B => n162, C => n6785, D => 
                           v_TEMP_VECTOR_7_port, Z => n161);
   U657 : AO7 port map( A => v_KEY_COL_OUT0_8_port, B => n121, C => n6781, Z =>
                           n152);
   U658 : AO7 port map( A => v_KEY_COL_OUT0_16_port, B => n80, C => n6783, Z =>
                           n111);
   U659 : AO7 port map( A => v_KEY_COL_OUT0_24_port, B => n21, C => n2501, Z =>
                           n61);
   U660 : AO7 port map( A => v_KEY_COL_OUT0_9_port, B => n121, C => n6781, Z =>
                           n146);
   U661 : AO7 port map( A => v_KEY_COL_OUT0_17_port, B => n80, C => n6783, Z =>
                           n105);
   U662 : AO7 port map( A => v_KEY_COL_OUT0_25_port, B => n21, C => n2501, Z =>
                           n52);
   U663 : AO7 port map( A => v_KEY_COL_OUT0_10_port, B => n121, C => n6781, Z 
                           => n142);
   U664 : AO7 port map( A => v_KEY_COL_OUT0_18_port, B => n80, C => n6783, Z =>
                           n101);
   U665 : AO7 port map( A => v_KEY_COL_OUT0_26_port, B => n21, C => n2501, Z =>
                           n47);
   U666 : AO7 port map( A => v_KEY_COL_OUT0_11_port, B => n121, C => n6781, Z 
                           => n138);
   U667 : AO7 port map( A => v_KEY_COL_OUT0_19_port, B => n80, C => n6783, Z =>
                           n97);
   U668 : AO7 port map( A => v_KEY_COL_OUT0_27_port, B => n21, C => n2501, Z =>
                           n42);
   U669 : AO7 port map( A => v_KEY_COL_OUT0_12_port, B => n121, C => n6781, Z 
                           => n134);
   U670 : AO7 port map( A => v_KEY_COL_OUT0_20_port, B => n80, C => n6783, Z =>
                           n93);
   U671 : AO7 port map( A => v_KEY_COL_OUT0_28_port, B => n21, C => n2501, Z =>
                           n37);
   U672 : AO7 port map( A => v_KEY_COL_OUT0_13_port, B => n121, C => n6781, Z 
                           => n130);
   U673 : AO7 port map( A => v_KEY_COL_OUT0_21_port, B => n80, C => n6783, Z =>
                           n89);
   U674 : AO7 port map( A => v_KEY_COL_OUT0_29_port, B => n21, C => n2501, Z =>
                           n32);
   U675 : AO7 port map( A => v_KEY_COL_OUT0_14_port, B => n121, C => n6781, Z 
                           => n126);
   U676 : AO7 port map( A => v_KEY_COL_OUT0_22_port, B => n80, C => n6783, Z =>
                           n85);
   U677 : AO7 port map( A => v_KEY_COL_OUT0_30_port, B => n21, C => n2501, Z =>
                           n27);
   U678 : AO7 port map( A => v_KEY_COL_OUT0_15_port, B => n121, C => n6781, Z 
                           => n120);
   U679 : AO7 port map( A => v_KEY_COL_OUT0_23_port, B => n80, C => n6783, Z =>
                           n79);
   U680 : AO7 port map( A => v_KEY_COL_OUT0_31_port, B => n21, C => n2501, Z =>
                           n20);
   U681 : AO3 port map( A => n2181, B => n114, C => n147, D => n148, Z => n6701
                           );
   U682 : AO2 port map( A => n151, B => v_KEY_COL_OUT0_8_port, C => 
                           v_TEMP_VECTOR_8_port, D => n152, Z => n147);
   U683 : AO2 port map( A => n117, B => v_TEMP_VECTOR_16_port, C => 
                           v_KEY32_IN_8_port, D => n118, Z => n148);
   U685 : AO3 port map( A => n2181, B => n73, C => n106, D => n107, Z => n6693)
                           ;
   U686 : AO2 port map( A => n110, B => v_KEY_COL_OUT0_16_port, C => 
                           v_TEMP_VECTOR_16_port, D => n111, Z => n106);
   U687 : AO2 port map( A => n76, B => v_TEMP_VECTOR_24_port, C => 
                           v_KEY32_IN_16_port, D => n77, Z => n107);
   U688 : AO3 port map( A => n13, B => n2181, C => n54, D => n55, Z => n6685);
   U689 : AO2 port map( A => n60, B => v_KEY_COL_OUT0_24_port, C => 
                           v_TEMP_VECTOR_24_port, D => n61, Z => n54);
   U690 : AO2 port map( A => v_TEMP_VECTOR_0_port, B => n17, C => 
                           v_KEY32_IN_24_port, D => n18, Z => n55);
   U691 : AO3 port map( A => n2205, B => n114, C => n143, D => n144, Z => n6700
                           );
   U692 : AO2 port map( A => n145, B => v_KEY_COL_OUT0_9_port, C => 
                           v_TEMP_VECTOR_9_port, D => n146, Z => n143);
   U693 : AO2 port map( A => n117, B => v_TEMP_VECTOR_17_port, C => 
                           v_KEY32_IN_9_port, D => n118, Z => n144);
   U694 : AO3 port map( A => n2205, B => n73, C => n102, D => n103, Z => n6692)
                           ;
   U695 : AO2 port map( A => n104, B => v_KEY_COL_OUT0_17_port, C => 
                           v_TEMP_VECTOR_17_port, D => n105, Z => n102);
   U696 : AO2 port map( A => n76, B => v_TEMP_VECTOR_25_port, C => 
                           v_KEY32_IN_17_port, D => n77, Z => n103);
   U697 : AO3 port map( A => n13, B => n2205, C => n49, D => n50, Z => n6684);
   U698 : AO2 port map( A => n51, B => v_KEY_COL_OUT0_25_port, C => 
                           v_TEMP_VECTOR_25_port, D => n52, Z => n49);
   U699 : AO2 port map( A => v_TEMP_VECTOR_1_port, B => n17, C => 
                           v_KEY32_IN_25_port, D => n18, Z => n50);
   U700 : AO3 port map( A => n2217, B => n114, C => n139, D => n140, Z => n6699
                           );
   U701 : AO2 port map( A => n141, B => v_KEY_COL_OUT0_10_port, C => 
                           v_TEMP_VECTOR_10_port, D => n142, Z => n139);
   U702 : AO2 port map( A => n117, B => v_TEMP_VECTOR_18_port, C => 
                           v_KEY32_IN_10_port, D => n118, Z => n140);
   U703 : AO3 port map( A => n2217, B => n73, C => n98, D => n99, Z => n6691);
   U704 : AO2 port map( A => n100, B => v_KEY_COL_OUT0_18_port, C => 
                           v_TEMP_VECTOR_18_port, D => n101, Z => n98);
   U705 : AO2 port map( A => n76, B => v_TEMP_VECTOR_26_port, C => 
                           v_KEY32_IN_18_port, D => n77, Z => n99);
   U706 : AO3 port map( A => n13, B => n2217, C => n44, D => n45, Z => n6683);
   U707 : AO2 port map( A => n46, B => v_KEY_COL_OUT0_26_port, C => 
                           v_TEMP_VECTOR_26_port, D => n47, Z => n44);
   U708 : AO2 port map( A => v_TEMP_VECTOR_2_port, B => n17, C => 
                           v_KEY32_IN_26_port, D => n18, Z => n45);
   U709 : AO3 port map( A => n2220, B => n114, C => n135, D => n136, Z => n6698
                           );
   U710 : AO2 port map( A => n137, B => v_KEY_COL_OUT0_11_port, C => 
                           v_TEMP_VECTOR_11_port, D => n138, Z => n135);
   U711 : AO2 port map( A => n117, B => v_TEMP_VECTOR_19_port, C => 
                           v_KEY32_IN_11_port, D => n118, Z => n136);
   U712 : AO3 port map( A => n2220, B => n73, C => n94, D => n95, Z => n6690);
   U713 : AO2 port map( A => n96, B => v_KEY_COL_OUT0_19_port, C => 
                           v_TEMP_VECTOR_19_port, D => n97, Z => n94);
   U714 : AO2 port map( A => n76, B => v_TEMP_VECTOR_27_port, C => 
                           v_KEY32_IN_19_port, D => n77, Z => n95);
   U715 : AO3 port map( A => n13, B => n2220, C => n39, D => n40, Z => n6682);
   U716 : AO2 port map( A => n41, B => v_KEY_COL_OUT0_27_port, C => 
                           v_TEMP_VECTOR_27_port, D => n42, Z => n39);
   U717 : AO2 port map( A => v_TEMP_VECTOR_3_port, B => n17, C => 
                           v_KEY32_IN_27_port, D => n18, Z => n40);
   U718 : AO3 port map( A => n2244, B => n114, C => n131, D => n132, Z => n6697
                           );
   U719 : AO2 port map( A => n133, B => v_KEY_COL_OUT0_12_port, C => 
                           v_TEMP_VECTOR_12_port, D => n134, Z => n131);
   U720 : AO2 port map( A => n117, B => v_TEMP_VECTOR_20_port, C => 
                           v_KEY32_IN_12_port, D => n118, Z => n132);
   U721 : AO3 port map( A => n2244, B => n73, C => n90, D => n91, Z => n6689);
   U722 : AO2 port map( A => n92, B => v_KEY_COL_OUT0_20_port, C => 
                           v_TEMP_VECTOR_20_port, D => n93, Z => n90);
   U723 : AO2 port map( A => n76, B => v_TEMP_VECTOR_28_port, C => 
                           v_KEY32_IN_20_port, D => n77, Z => n91);
   U724 : AO3 port map( A => n13, B => n2244, C => n34, D => n35, Z => n6681);
   U725 : AO2 port map( A => n36, B => v_KEY_COL_OUT0_28_port, C => 
                           v_TEMP_VECTOR_28_port, D => n37, Z => n34);
   U726 : AO2 port map( A => v_TEMP_VECTOR_4_port, B => n17, C => 
                           v_KEY32_IN_28_port, D => n18, Z => n35);
   U727 : AO3 port map( A => n2233, B => n114, C => n127, D => n128, Z => n6696
                           );
   U729 : AO2 port map( A => n129, B => v_KEY_COL_OUT0_13_port, C => 
                           v_TEMP_VECTOR_13_port, D => n130, Z => n127);
   U730 : AO2 port map( A => n117, B => v_TEMP_VECTOR_21_port, C => 
                           v_KEY32_IN_13_port, D => n118, Z => n128);
   U731 : AO3 port map( A => n2233, B => n73, C => n86, D => n87, Z => n6688);
   U732 : AO2 port map( A => n88, B => v_KEY_COL_OUT0_21_port, C => 
                           v_TEMP_VECTOR_21_port, D => n89, Z => n86);
   U733 : AO2 port map( A => n76, B => v_TEMP_VECTOR_29_port, C => 
                           v_KEY32_IN_21_port, D => n77, Z => n87);
   U734 : AO3 port map( A => n13, B => n2233, C => n29, D => n30, Z => n6680);
   U735 : AO2 port map( A => n31, B => v_KEY_COL_OUT0_29_port, C => 
                           v_TEMP_VECTOR_29_port, D => n32, Z => n29);
   U736 : AO2 port map( A => v_TEMP_VECTOR_5_port, B => n17, C => 
                           v_KEY32_IN_29_port, D => n18, Z => n30);
   U737 : AO3 port map( A => n2183, B => n114, C => n123, D => n124, Z => n6695
                           );
   U738 : AO2 port map( A => n125, B => v_KEY_COL_OUT0_14_port, C => 
                           v_TEMP_VECTOR_14_port, D => n126, Z => n123);
   U739 : AO2 port map( A => n117, B => v_TEMP_VECTOR_22_port, C => 
                           v_KEY32_IN_14_port, D => n118, Z => n124);
   U740 : AO3 port map( A => n2183, B => n73, C => n82, D => n83, Z => n6687);
   U741 : AO2 port map( A => n84, B => v_KEY_COL_OUT0_22_port, C => 
                           v_TEMP_VECTOR_22_port, D => n85, Z => n82);
   U742 : AO2 port map( A => n76, B => v_TEMP_VECTOR_30_port, C => 
                           v_KEY32_IN_22_port, D => n77, Z => n83);
   U743 : AO3 port map( A => n13, B => n2183, C => n24, D => n25, Z => n6679);
   U744 : AO2 port map( A => n26, B => v_KEY_COL_OUT0_30_port, C => 
                           v_TEMP_VECTOR_30_port, D => n27, Z => n24);
   U745 : AO2 port map( A => v_TEMP_VECTOR_6_port, B => n17, C => 
                           v_KEY32_IN_30_port, D => n18, Z => n25);
   U746 : AO3 port map( A => n2240, B => n114, C => n115, D => n116, Z => n6694
                           );
   U747 : AO2 port map( A => n119, B => v_KEY_COL_OUT0_15_port, C => 
                           v_TEMP_VECTOR_15_port, D => n120, Z => n115);
   U748 : AO2 port map( A => n117, B => v_TEMP_VECTOR_23_port, C => 
                           v_KEY32_IN_15_port, D => n118, Z => n116);
   U749 : AO3 port map( A => n2240, B => n73, C => n74, D => n75, Z => n6686);
   U750 : AO2 port map( A => n78, B => v_KEY_COL_OUT0_23_port, C => 
                           v_TEMP_VECTOR_23_port, D => n79, Z => n74);
   U751 : AO2 port map( A => n76, B => v_TEMP_VECTOR_31_port, C => 
                           v_KEY32_IN_23_port, D => n77, Z => n75);
   U752 : AO3 port map( A => n13, B => n2240, C => n15, D => n16, Z => n6678);
   U753 : AO2 port map( A => n19, B => v_KEY_COL_OUT0_31_port, C => 
                           v_TEMP_VECTOR_31_port, D => n20, Z => n15);
   U754 : AO2 port map( A => v_TEMP_VECTOR_7_port, B => n17, C => 
                           v_KEY32_IN_31_port, D => n18, Z => n16);
   U755 : AO2 port map( A => v_TEMP_VECTOR_24_port, B => n112, C => 
                           v_TEMP_VECTOR_16_port, D => n153, Z => n2296);
   U756 : AO2 port map( A => v_TEMP_VECTOR_8_port, B => n1876, C => 
                           v_TEMP_VECTOR_0_port, D => n2281, Z => n2295);
   U757 : AO2 port map( A => v_KEY32_IN_8_port, B => n1543, C => 
                           v_TEMP_VECTOR_8_port, D => n1499, Z => n2446);
   U758 : AO2 port map( A => v_KEY32_IN_16_port, B => n1543, C => 
                           v_TEMP_VECTOR_16_port, D => n1499, Z => n2454);
   U759 : AO2 port map( A => v_KEY32_IN_24_port, B => n1543, C => 
                           v_TEMP_VECTOR_24_port, D => n1499, Z => n2462);
   U760 : AO2 port map( A => v_KEY32_IN_9_port, B => n1543, C => 
                           v_TEMP_VECTOR_9_port, D => n1499, Z => n2447);
   U761 : AO2 port map( A => v_KEY32_IN_17_port, B => n1543, C => 
                           v_TEMP_VECTOR_17_port, D => n1499, Z => n2455);
   U762 : AO2 port map( A => v_KEY32_IN_25_port, B => n1543, C => 
                           v_TEMP_VECTOR_25_port, D => n1499, Z => n2463);
   U763 : AO2 port map( A => v_KEY32_IN_10_port, B => n1543, C => 
                           v_TEMP_VECTOR_10_port, D => n1499, Z => n2448);
   U764 : AO2 port map( A => v_KEY32_IN_18_port, B => n1543, C => 
                           v_TEMP_VECTOR_18_port, D => n1499, Z => n2456);
   U765 : AO2 port map( A => v_KEY32_IN_26_port, B => n1543, C => 
                           v_TEMP_VECTOR_26_port, D => n1499, Z => n2464);
   U766 : AO2 port map( A => v_KEY32_IN_11_port, B => n1543, C => 
                           v_TEMP_VECTOR_11_port, D => n1499, Z => n2449);
   U767 : AO2 port map( A => v_KEY32_IN_19_port, B => n1543, C => 
                           v_TEMP_VECTOR_19_port, D => n1499, Z => n2457);
   U768 : AO2 port map( A => v_KEY32_IN_27_port, B => n1543, C => 
                           v_TEMP_VECTOR_27_port, D => n1499, Z => n2465);
   U769 : AO2 port map( A => v_KEY32_IN_12_port, B => n1543, C => 
                           v_TEMP_VECTOR_12_port, D => n1499, Z => n2450);
   U770 : AO2 port map( A => v_KEY32_IN_20_port, B => n1543, C => 
                           v_TEMP_VECTOR_20_port, D => n1499, Z => n2458);
   U771 : AO2 port map( A => v_KEY32_IN_28_port, B => n1543, C => 
                           v_TEMP_VECTOR_28_port, D => n1499, Z => n2466);
   U773 : AO2 port map( A => v_KEY32_IN_4_port, B => n1543, C => 
                           v_TEMP_VECTOR_4_port, D => n1499, Z => n2442);
   U774 : AO2 port map( A => v_KEY32_IN_13_port, B => n1543, C => 
                           v_TEMP_VECTOR_13_port, D => n1499, Z => n2451);
   U775 : AO2 port map( A => v_KEY32_IN_21_port, B => n1543, C => 
                           v_TEMP_VECTOR_21_port, D => n1499, Z => n2459);
   U776 : AO2 port map( A => v_KEY32_IN_29_port, B => n1543, C => 
                           v_TEMP_VECTOR_29_port, D => n1499, Z => n2467);
   U777 : AO2 port map( A => v_KEY32_IN_5_port, B => n1543, C => 
                           v_TEMP_VECTOR_5_port, D => n1499, Z => n2443);
   U778 : AO2 port map( A => v_KEY32_IN_14_port, B => n1543, C => 
                           v_TEMP_VECTOR_14_port, D => n1499, Z => n2452);
   U779 : AO2 port map( A => v_KEY32_IN_22_port, B => n1543, C => 
                           v_TEMP_VECTOR_22_port, D => n1499, Z => n2460);
   U780 : AO2 port map( A => v_KEY32_IN_30_port, B => n1543, C => 
                           v_TEMP_VECTOR_30_port, D => n1499, Z => n2468);
   U781 : AO2 port map( A => v_KEY32_IN_6_port, B => n1543, C => 
                           v_TEMP_VECTOR_6_port, D => n1499, Z => n2444);
   U782 : AO2 port map( A => v_KEY32_IN_15_port, B => n1543, C => 
                           v_TEMP_VECTOR_15_port, D => n1499, Z => n2453);
   U783 : AO2 port map( A => v_KEY32_IN_23_port, B => n1543, C => 
                           v_TEMP_VECTOR_23_port, D => n1499, Z => n2461);
   U784 : AO2 port map( A => v_KEY32_IN_31_port, B => n1543, C => 
                           v_TEMP_VECTOR_31_port, D => n1499, Z => n2469);
   U785 : AO2 port map( A => v_KEY32_IN_7_port, B => n1543, C => 
                           v_TEMP_VECTOR_7_port, D => n1499, Z => n2445);
   U786 : AO4 port map( A => n2548, B => n378, C => n375, D => n2390, Z => 
                           n5117);
   U787 : AO4 port map( A => n2549, B => n383, C => n2446, D => n2389, Z => 
                           n5118);
   U788 : AO4 port map( A => n2546, B => n384, C => n2446, D => n2388, Z => 
                           n5119);
   U789 : AO4 port map( A => n2547, B => n385, C => n2446, D => n2387, Z => 
                           n5120);
   U790 : AO4 port map( A => n2544, B => n386, C => n375, D => n2386, Z => 
                           n5121);
   U791 : AO4 port map( A => n2545, B => n387, C => n2446, D => n2385, Z => 
                           n5122);
   U792 : AO4 port map( A => n2542, B => n388, C => n2446, D => n2384, Z => 
                           n5123);
   U793 : AO4 port map( A => n2543, B => n389, C => n2446, D => n2383, Z => 
                           n5124);
   U794 : AO4 port map( A => n2612, B => n378, C => n2454, D => n2390, Z => 
                           n5629);
   U795 : AO4 port map( A => n2613, B => n383, C => n374, D => n2389, Z => 
                           n5630);
   U796 : AO4 port map( A => n2610, B => n384, C => n2454, D => n2388, Z => 
                           n5631);
   U797 : AO4 port map( A => n2611, B => n385, C => n2454, D => n2387, Z => 
                           n5632);
   U798 : AO4 port map( A => n2608, B => n386, C => n374, D => n2386, Z => 
                           n5633);
   U799 : AO4 port map( A => n2609, B => n387, C => n2454, D => n2385, Z => 
                           n5634);
   U800 : AO4 port map( A => n2606, B => n388, C => n2454, D => n2384, Z => 
                           n5635);
   U801 : AO4 port map( A => n2607, B => n389, C => n2454, D => n2383, Z => 
                           n5636);
   U802 : AO4 port map( A => n2676, B => n378, C => n2462, D => n2390, Z => 
                           n6141);
   U803 : AO4 port map( A => n2677, B => n383, C => n351, D => n2389, Z => 
                           n6142);
   U804 : AO4 port map( A => n2674, B => n384, C => n2462, D => n2388, Z => 
                           n6143);
   U805 : AO4 port map( A => n2675, B => n385, C => n2462, D => n2387, Z => 
                           n6144);
   U806 : AO4 port map( A => n2672, B => n386, C => n351, D => n2386, Z => 
                           n6145);
   U807 : AO4 port map( A => n2673, B => n387, C => n2462, D => n2385, Z => 
                           n6146);
   U808 : AO4 port map( A => n2670, B => n388, C => n2462, D => n2384, Z => 
                           n6147);
   U809 : AO4 port map( A => n2671, B => n389, C => n2462, D => n2383, Z => 
                           n6148);
   U810 : AO4 port map( A => n2804, B => n378, C => n373, D => n2390, Z => 
                           n5181);
   U811 : AO4 port map( A => n2805, B => n383, C => n2447, D => n2389, Z => 
                           n5182);
   U812 : AO4 port map( A => n2802, B => n384, C => n2447, D => n2388, Z => 
                           n5183);
   U813 : AO4 port map( A => n2803, B => n385, C => n2447, D => n2387, Z => 
                           n5184);
   U814 : AO4 port map( A => n2800, B => n386, C => n373, D => n2386, Z => 
                           n5185);
   U815 : AO4 port map( A => n2801, B => n387, C => n2447, D => n2385, Z => 
                           n5186);
   U817 : AO4 port map( A => n2798, B => n388, C => n2447, D => n2384, Z => 
                           n5187);
   U818 : AO4 port map( A => n2799, B => n389, C => n2447, D => n2383, Z => 
                           n5188);
   U819 : AO4 port map( A => n2868, B => n378, C => n372, D => n2390, Z => 
                           n5693);
   U820 : AO4 port map( A => n2869, B => n383, C => n2455, D => n2389, Z => 
                           n5694);
   U821 : AO4 port map( A => n2866, B => n384, C => n2455, D => n2388, Z => 
                           n5695);
   U822 : AO4 port map( A => n2867, B => n385, C => n2455, D => n2387, Z => 
                           n5696);
   U823 : AO4 port map( A => n2864, B => n386, C => n372, D => n2386, Z => 
                           n5697);
   U824 : AO4 port map( A => n2865, B => n387, C => n2455, D => n2385, Z => 
                           n5698);
   U825 : AO4 port map( A => n2862, B => n388, C => n2455, D => n2384, Z => 
                           n5699);
   U826 : AO4 port map( A => n2863, B => n389, C => n2455, D => n2383, Z => 
                           n5700);
   U827 : AO4 port map( A => n2932, B => n378, C => n350, D => n2390, Z => 
                           n6205);
   U828 : AO4 port map( A => n2933, B => n383, C => n2463, D => n2389, Z => 
                           n6206);
   U829 : AO4 port map( A => n2930, B => n384, C => n2463, D => n2388, Z => 
                           n6207);
   U830 : AO4 port map( A => n2931, B => n385, C => n2463, D => n2387, Z => 
                           n6208);
   U831 : AO4 port map( A => n2928, B => n386, C => n350, D => n2386, Z => 
                           n6209);
   U832 : AO4 port map( A => n2929, B => n387, C => n2463, D => n2385, Z => 
                           n6210);
   U833 : AO4 port map( A => n2926, B => n388, C => n2463, D => n2384, Z => 
                           n6211);
   U834 : AO4 port map( A => n2927, B => n389, C => n2463, D => n2383, Z => 
                           n6212);
   U835 : AO4 port map( A => n3060, B => n378, C => n2448, D => n2390, Z => 
                           n5245);
   U836 : AO4 port map( A => n3061, B => n383, C => n2448, D => n2389, Z => 
                           n5246);
   U837 : AO4 port map( A => n3058, B => n384, C => n2448, D => n2388, Z => 
                           n5247);
   U838 : AO4 port map( A => n3059, B => n385, C => n2448, D => n2387, Z => 
                           n5248);
   U839 : AO4 port map( A => n3056, B => n386, C => n2448, D => n2386, Z => 
                           n5249);
   U840 : AO4 port map( A => n3057, B => n387, C => n2448, D => n2385, Z => 
                           n5250);
   U841 : AO4 port map( A => n3054, B => n388, C => n2448, D => n2384, Z => 
                           n5251);
   U842 : AO4 port map( A => n3055, B => n389, C => n2448, D => n2383, Z => 
                           n5252);
   U843 : AO4 port map( A => n3124, B => n378, C => n349, D => n2390, Z => 
                           n5757);
   U844 : AO4 port map( A => n3125, B => n383, C => n2456, D => n2389, Z => 
                           n5758);
   U845 : AO4 port map( A => n3122, B => n384, C => n2456, D => n2388, Z => 
                           n5759);
   U846 : AO4 port map( A => n3123, B => n385, C => n2456, D => n2387, Z => 
                           n5760);
   U847 : AO4 port map( A => n3120, B => n386, C => n349, D => n2386, Z => 
                           n5761);
   U848 : AO4 port map( A => n3121, B => n387, C => n2456, D => n2385, Z => 
                           n5762);
   U849 : AO4 port map( A => n3118, B => n388, C => n2456, D => n2384, Z => 
                           n5763);
   U850 : AO4 port map( A => n3119, B => n389, C => n2456, D => n2383, Z => 
                           n5764);
   U851 : AO4 port map( A => n3188, B => n378, C => n2464, D => n2390, Z => 
                           n6269);
   U852 : AO4 port map( A => n3189, B => n383, C => n2464, D => n2389, Z => 
                           n6270);
   U853 : AO4 port map( A => n3186, B => n384, C => n2464, D => n2388, Z => 
                           n6271);
   U854 : AO4 port map( A => n3187, B => n385, C => n2464, D => n2387, Z => 
                           n6272);
   U855 : AO4 port map( A => n3184, B => n386, C => n2464, D => n2386, Z => 
                           n6273);
   U856 : AO4 port map( A => n3185, B => n387, C => n2464, D => n2385, Z => 
                           n6274);
   U857 : AO4 port map( A => n3182, B => n388, C => n2464, D => n2384, Z => 
                           n6275);
   U858 : AO4 port map( A => n3183, B => n389, C => n2464, D => n2383, Z => 
                           n6276);
   U859 : AO4 port map( A => n3316, B => n378, C => n366, D => n2390, Z => 
                           n5309);
   U861 : AO4 port map( A => n3317, B => n383, C => n2449, D => n2389, Z => 
                           n5310);
   U862 : AO4 port map( A => n3314, B => n384, C => n2449, D => n2388, Z => 
                           n5311);
   U863 : AO4 port map( A => n3315, B => n385, C => n2449, D => n2387, Z => 
                           n5312);
   U864 : AO4 port map( A => n3312, B => n386, C => n366, D => n2386, Z => 
                           n5313);
   U865 : AO4 port map( A => n3313, B => n387, C => n2449, D => n2385, Z => 
                           n5314);
   U866 : AO4 port map( A => n3310, B => n388, C => n2449, D => n2384, Z => 
                           n5315);
   U867 : AO4 port map( A => n3311, B => n389, C => n2449, D => n2383, Z => 
                           n5316);
   U868 : AO4 port map( A => n3380, B => n378, C => n347, D => n2390, Z => 
                           n5821);
   U869 : AO4 port map( A => n3381, B => n383, C => n2457, D => n2389, Z => 
                           n5822);
   U870 : AO4 port map( A => n3378, B => n384, C => n2457, D => n2388, Z => 
                           n5823);
   U871 : AO4 port map( A => n3379, B => n385, C => n2457, D => n2387, Z => 
                           n5824);
   U872 : AO4 port map( A => n3376, B => n386, C => n347, D => n2386, Z => 
                           n5825);
   U873 : AO4 port map( A => n3377, B => n387, C => n2457, D => n2385, Z => 
                           n5826);
   U874 : AO4 port map( A => n3374, B => n388, C => n2457, D => n2384, Z => 
                           n5827);
   U875 : AO4 port map( A => n3375, B => n389, C => n2457, D => n2383, Z => 
                           n5828);
   U876 : AO4 port map( A => n3444, B => n378, C => n2465, D => n2390, Z => 
                           n6333);
   U877 : AO4 port map( A => n3445, B => n383, C => n335, D => n2389, Z => 
                           n6334);
   U878 : AO4 port map( A => n3442, B => n384, C => n2465, D => n2388, Z => 
                           n6335);
   U879 : AO4 port map( A => n3443, B => n385, C => n2465, D => n2387, Z => 
                           n6336);
   U880 : AO4 port map( A => n3440, B => n386, C => n335, D => n2386, Z => 
                           n6337);
   U881 : AO4 port map( A => n3441, B => n387, C => n2465, D => n2385, Z => 
                           n6338);
   U882 : AO4 port map( A => n3438, B => n388, C => n2465, D => n2384, Z => 
                           n6339);
   U883 : AO4 port map( A => n3439, B => n389, C => n2465, D => n2383, Z => 
                           n6340);
   U884 : AO4 port map( A => n3572, B => n378, C => n2450, D => n2390, Z => 
                           n5373);
   U885 : AO4 port map( A => n3573, B => n383, C => n365, D => n2389, Z => 
                           n5374);
   U886 : AO4 port map( A => n3570, B => n384, C => n2450, D => n2388, Z => 
                           n5375);
   U887 : AO4 port map( A => n3571, B => n385, C => n2450, D => n2387, Z => 
                           n5376);
   U888 : AO4 port map( A => n3568, B => n386, C => n365, D => n2386, Z => 
                           n5377);
   U889 : AO4 port map( A => n3569, B => n387, C => n2450, D => n2385, Z => 
                           n5378);
   U890 : AO4 port map( A => n3566, B => n388, C => n2450, D => n2384, Z => 
                           n5379);
   U891 : AO4 port map( A => n3567, B => n389, C => n2450, D => n2383, Z => 
                           n5380);
   U892 : AO4 port map( A => n3636, B => n378, C => n325, D => n2390, Z => 
                           n5885);
   U893 : AO4 port map( A => n3637, B => n383, C => n2458, D => n2389, Z => 
                           n5886);
   U894 : AO4 port map( A => n3634, B => n384, C => n2458, D => n2388, Z => 
                           n5887);
   U895 : AO4 port map( A => n3635, B => n385, C => n2458, D => n2387, Z => 
                           n5888);
   U896 : AO4 port map( A => n3632, B => n386, C => n325, D => n2386, Z => 
                           n5889);
   U897 : AO4 port map( A => n3633, B => n387, C => n2458, D => n2385, Z => 
                           n5890);
   U898 : AO4 port map( A => n3630, B => n388, C => n2458, D => n2384, Z => 
                           n5891);
   U899 : AO4 port map( A => n3631, B => n389, C => n2458, D => n2383, Z => 
                           n5892);
   U900 : AO4 port map( A => n3700, B => n378, C => n314, D => n2390, Z => 
                           n6397);
   U901 : AO4 port map( A => n3701, B => n383, C => n2466, D => n2389, Z => 
                           n6398);
   U902 : AO4 port map( A => n3698, B => n384, C => n2466, D => n2388, Z => 
                           n6399);
   U903 : AO4 port map( A => n3699, B => n385, C => n2466, D => n2387, Z => 
                           n6400);
   U905 : AO4 port map( A => n3696, B => n386, C => n314, D => n2386, Z => 
                           n6401);
   U906 : AO4 port map( A => n3697, B => n387, C => n2466, D => n2385, Z => 
                           n6402);
   U907 : AO4 port map( A => n3694, B => n388, C => n2466, D => n2384, Z => 
                           n6403);
   U908 : AO4 port map( A => n3695, B => n389, C => n2466, D => n2383, Z => 
                           n6404);
   U909 : AO4 port map( A => n3764, B => n378, C => n364, D => n2390, Z => 
                           n4861);
   U910 : AO4 port map( A => n3765, B => n383, C => n2442, D => n2389, Z => 
                           n4862);
   U911 : AO4 port map( A => n3762, B => n384, C => n2442, D => n2388, Z => 
                           n4863);
   U912 : AO4 port map( A => n3763, B => n385, C => n2442, D => n2387, Z => 
                           n4864);
   U913 : AO4 port map( A => n3760, B => n386, C => n364, D => n2386, Z => 
                           n4865);
   U914 : AO4 port map( A => n3761, B => n387, C => n2442, D => n2385, Z => 
                           n4866);
   U915 : AO4 port map( A => n3758, B => n388, C => n2442, D => n2384, Z => 
                           n4867);
   U916 : AO4 port map( A => n3759, B => n389, C => n2442, D => n2383, Z => 
                           n4868);
   U917 : AO4 port map( A => n3828, B => n378, C => n363, D => n2390, Z => 
                           n5437);
   U918 : AO4 port map( A => n3829, B => n383, C => n2451, D => n2389, Z => 
                           n5438);
   U919 : AO4 port map( A => n3826, B => n384, C => n2451, D => n2388, Z => 
                           n5439);
   U920 : AO4 port map( A => n3827, B => n385, C => n2451, D => n2387, Z => 
                           n5440);
   U921 : AO4 port map( A => n3824, B => n386, C => n363, D => n2386, Z => 
                           n5441);
   U922 : AO4 port map( A => n3825, B => n387, C => n2451, D => n2385, Z => 
                           n5442);
   U923 : AO4 port map( A => n3822, B => n388, C => n2451, D => n2384, Z => 
                           n5443);
   U924 : AO4 port map( A => n3823, B => n389, C => n2451, D => n2383, Z => 
                           n5444);
   U925 : AO4 port map( A => n3892, B => n378, C => n2459, D => n2390, Z => 
                           n5949);
   U926 : AO4 port map( A => n3893, B => n383, C => n2459, D => n2389, Z => 
                           n5950);
   U927 : AO4 port map( A => n3890, B => n384, C => n2459, D => n2388, Z => 
                           n5951);
   U928 : AO4 port map( A => n3891, B => n385, C => n2459, D => n2387, Z => 
                           n5952);
   U929 : AO4 port map( A => n3888, B => n386, C => n2459, D => n2386, Z => 
                           n5953);
   U930 : AO4 port map( A => n3889, B => n387, C => n2459, D => n2385, Z => 
                           n5954);
   U931 : AO4 port map( A => n3886, B => n388, C => n2459, D => n2384, Z => 
                           n5955);
   U932 : AO4 port map( A => n3887, B => n389, C => n2459, D => n2383, Z => 
                           n5956);
   U933 : AO4 port map( A => n3956, B => n378, C => n301, D => n2390, Z => 
                           n6461);
   U934 : AO4 port map( A => n3957, B => n383, C => n2467, D => n2389, Z => 
                           n6462);
   U935 : AO4 port map( A => n3954, B => n384, C => n2467, D => n2388, Z => 
                           n6463);
   U936 : AO4 port map( A => n3955, B => n385, C => n2467, D => n2387, Z => 
                           n6464);
   U937 : AO4 port map( A => n3952, B => n386, C => n301, D => n2386, Z => 
                           n6465);
   U938 : AO4 port map( A => n3953, B => n387, C => n2467, D => n2385, Z => 
                           n6466);
   U939 : AO4 port map( A => n3950, B => n388, C => n2467, D => n2384, Z => 
                           n6467);
   U940 : AO4 port map( A => n3951, B => n389, C => n2467, D => n2383, Z => 
                           n6468);
   U941 : AO4 port map( A => n4020, B => n378, C => n2443, D => n2390, Z => 
                           n4925);
   U942 : AO4 port map( A => n4021, B => n383, C => n2443, D => n2389, Z => 
                           n4926);
   U943 : AO4 port map( A => n4018, B => n384, C => n2443, D => n2388, Z => 
                           n4927);
   U944 : AO4 port map( A => n4019, B => n385, C => n2443, D => n2387, Z => 
                           n4928);
   U945 : AO4 port map( A => n4016, B => n386, C => n2443, D => n2386, Z => 
                           n4929);
   U946 : AO4 port map( A => n4017, B => n387, C => n2443, D => n2385, Z => 
                           n4930);
   U947 : AO4 port map( A => n4014, B => n388, C => n2443, D => n2384, Z => 
                           n4931);
   U949 : AO4 port map( A => n4015, B => n389, C => n2443, D => n2383, Z => 
                           n4932);
   U950 : AO4 port map( A => n4084, B => n378, C => n361, D => n2390, Z => 
                           n5501);
   U951 : AO4 port map( A => n4085, B => n383, C => n2452, D => n2389, Z => 
                           n5502);
   U952 : AO4 port map( A => n4082, B => n384, C => n2452, D => n2388, Z => 
                           n5503);
   U953 : AO4 port map( A => n4083, B => n385, C => n2452, D => n2387, Z => 
                           n5504);
   U954 : AO4 port map( A => n4080, B => n386, C => n361, D => n2386, Z => 
                           n5505);
   U955 : AO4 port map( A => n4081, B => n387, C => n2452, D => n2385, Z => 
                           n5506);
   U956 : AO4 port map( A => n4078, B => n388, C => n2452, D => n2384, Z => 
                           n5507);
   U957 : AO4 port map( A => n4079, B => n389, C => n2452, D => n2383, Z => 
                           n5508);
   U958 : AO4 port map( A => n4148, B => n378, C => n2460, D => n2390, Z => 
                           n6013);
   U959 : AO4 port map( A => n4149, B => n383, C => n293, D => n2389, Z => 
                           n6014);
   U960 : AO4 port map( A => n4146, B => n384, C => n2460, D => n2388, Z => 
                           n6015);
   U961 : AO4 port map( A => n4147, B => n385, C => n2460, D => n2387, Z => 
                           n6016);
   U962 : AO4 port map( A => n4144, B => n386, C => n293, D => n2386, Z => 
                           n6017);
   U963 : AO4 port map( A => n4145, B => n387, C => n2460, D => n2385, Z => 
                           n6018);
   U964 : AO4 port map( A => n4142, B => n388, C => n2460, D => n2384, Z => 
                           n6019);
   U965 : AO4 port map( A => n4143, B => n389, C => n2460, D => n2383, Z => 
                           n6020);
   U966 : AO4 port map( A => n4212, B => n378, C => n286, D => n2390, Z => 
                           n6525);
   U967 : AO4 port map( A => n4213, B => n383, C => n2468, D => n2389, Z => 
                           n6526);
   U968 : AO4 port map( A => n4210, B => n384, C => n2468, D => n2388, Z => 
                           n6527);
   U969 : AO4 port map( A => n4211, B => n385, C => n2468, D => n2387, Z => 
                           n6528);
   U970 : AO4 port map( A => n4208, B => n386, C => n286, D => n2386, Z => 
                           n6529);
   U971 : AO4 port map( A => n4209, B => n387, C => n2468, D => n2385, Z => 
                           n6530);
   U972 : AO4 port map( A => n4206, B => n388, C => n2468, D => n2384, Z => 
                           n6531);
   U973 : AO4 port map( A => n4207, B => n389, C => n2468, D => n2383, Z => 
                           n6532);
   U974 : AO4 port map( A => n4276, B => n378, C => n2444, D => n2390, Z => 
                           n4989);
   U975 : AO4 port map( A => n4277, B => n383, C => n360, D => n2389, Z => 
                           n4990);
   U976 : AO4 port map( A => n4274, B => n384, C => n2444, D => n2388, Z => 
                           n4991);
   U977 : AO4 port map( A => n4275, B => n385, C => n2444, D => n2387, Z => 
                           n4992);
   U978 : AO4 port map( A => n4272, B => n386, C => n360, D => n2386, Z => 
                           n4993);
   U979 : AO4 port map( A => n4273, B => n387, C => n2444, D => n2385, Z => 
                           n4994);
   U980 : AO4 port map( A => n4270, B => n388, C => n2444, D => n2384, Z => 
                           n4995);
   U981 : AO4 port map( A => n4271, B => n389, C => n2444, D => n2383, Z => 
                           n4996);
   U982 : AO4 port map( A => n4340, B => n378, C => n359, D => n2390, Z => 
                           n5565);
   U983 : AO4 port map( A => n4341, B => n383, C => n2453, D => n2389, Z => 
                           n5566);
   U984 : AO4 port map( A => n4338, B => n384, C => n2453, D => n2388, Z => 
                           n5567);
   U985 : AO4 port map( A => n4339, B => n385, C => n2453, D => n2387, Z => 
                           n5568);
   U986 : AO4 port map( A => n4336, B => n386, C => n359, D => n2386, Z => 
                           n5569);
   U987 : AO4 port map( A => n4337, B => n387, C => n2453, D => n2385, Z => 
                           n5570);
   U988 : AO4 port map( A => n4334, B => n388, C => n2453, D => n2384, Z => 
                           n5571);
   U989 : AO4 port map( A => n4335, B => n389, C => n2453, D => n2383, Z => 
                           n5572);
   U990 : AO4 port map( A => n4404, B => n378, C => n284, D => n2390, Z => 
                           n6077);
   U991 : AO4 port map( A => n4405, B => n383, C => n2461, D => n2389, Z => 
                           n6078);
   U993 : AO4 port map( A => n4402, B => n384, C => n2461, D => n2388, Z => 
                           n6079);
   U994 : AO4 port map( A => n4403, B => n385, C => n2461, D => n2387, Z => 
                           n6080);
   U995 : AO4 port map( A => n4400, B => n386, C => n284, D => n2386, Z => 
                           n6081);
   U996 : AO4 port map( A => n4401, B => n387, C => n2461, D => n2385, Z => 
                           n6082);
   U997 : AO4 port map( A => n4398, B => n388, C => n2461, D => n2384, Z => 
                           n6083);
   U998 : AO4 port map( A => n4399, B => n389, C => n2461, D => n2383, Z => 
                           n6084);
   U999 : AO4 port map( A => n4468, B => n378, C => n2469, D => n2390, Z => 
                           n6589);
   U1000 : AO4 port map( A => n4469, B => n383, C => n2469, D => n2389, Z => 
                           n6590);
   U1001 : AO4 port map( A => n4466, B => n384, C => n2469, D => n2388, Z => 
                           n6591);
   U1002 : AO4 port map( A => n4467, B => n385, C => n2469, D => n2387, Z => 
                           n6592);
   U1003 : AO4 port map( A => n4464, B => n386, C => n2469, D => n2386, Z => 
                           n6593);
   U1004 : AO4 port map( A => n4465, B => n387, C => n2469, D => n2385, Z => 
                           n6594);
   U1005 : AO4 port map( A => n4462, B => n388, C => n2469, D => n2384, Z => 
                           n6595);
   U1006 : AO4 port map( A => n4463, B => n389, C => n2469, D => n2383, Z => 
                           n6596);
   U1007 : AO4 port map( A => n4532, B => n378, C => n354, D => n2390, Z => 
                           n5053);
   U1008 : AO4 port map( A => n4533, B => n383, C => n2445, D => n2389, Z => 
                           n5054);
   U1009 : AO4 port map( A => n4530, B => n384, C => n2445, D => n2388, Z => 
                           n5055);
   U1010 : AO4 port map( A => n4531, B => n385, C => n2445, D => n2387, Z => 
                           n5056);
   U1011 : AO4 port map( A => n4528, B => n386, C => n354, D => n2386, Z => 
                           n5057);
   U1012 : AO4 port map( A => n4529, B => n387, C => n2445, D => n2385, Z => 
                           n5058);
   U1013 : AO4 port map( A => n4526, B => n388, C => n2445, D => n2384, Z => 
                           n5059);
   U1014 : AO4 port map( A => n4527, B => n389, C => n2445, D => n2383, Z => 
                           n5060);
   U1015 : AO2 port map( A => v_KEY32_IN_0_port, B => n1543, C => 
                           v_TEMP_VECTOR_0_port, D => n1499, Z => n2309);
   U1016 : AO2 port map( A => v_KEY32_IN_1_port, B => n1543, C => 
                           v_TEMP_VECTOR_1_port, D => n1499, Z => n2439);
   U1017 : AO2 port map( A => v_KEY32_IN_2_port, B => n1543, C => 
                           v_TEMP_VECTOR_2_port, D => n1499, Z => n2440);
   U1018 : AO2 port map( A => v_KEY32_IN_3_port, B => n1543, C => 
                           v_TEMP_VECTOR_3_port, D => n1499, Z => n2441);
   U1019 : AO4 port map( A => n2556, B => n390, C => n375, D => n2382, Z => 
                           n5125);
   U1020 : AO4 port map( A => n2557, B => n399, C => n2446, D => n2381, Z => 
                           n5126);
   U1021 : AO4 port map( A => n2554, B => n400, C => n375, D => n2380, Z => 
                           n5127);
   U1022 : AO4 port map( A => n2555, B => n401, C => n2446, D => n2379, Z => 
                           n5128);
   U1023 : AO4 port map( A => n2552, B => n402, C => n375, D => n2378, Z => 
                           n5129);
   U1024 : AO4 port map( A => n2553, B => n403, C => n2446, D => n2377, Z => 
                           n5130);
   U1025 : AO4 port map( A => n2550, B => n404, C => n375, D => n2376, Z => 
                           n5131);
   U1026 : AO4 port map( A => n2551, B => n405, C => n2446, D => n2375, Z => 
                           n5132);
   U1027 : AO4 port map( A => n2564, B => n406, C => n375, D => n2374, Z => 
                           n5133);
   U1028 : AO4 port map( A => n2565, B => n411, C => n2446, D => n2373, Z => 
                           n5134);
   U1029 : AO4 port map( A => n2562, B => n412, C => n2446, D => n2372, Z => 
                           n5135);
   U1030 : AO4 port map( A => n2563, B => n413, C => n2446, D => n2371, Z => 
                           n5136);
   U1031 : AO4 port map( A => n2560, B => n414, C => n2446, D => n2370, Z => 
                           n5137);
   U1032 : AO4 port map( A => n2561, B => n415, C => n2446, D => n2369, Z => 
                           n5138);
   U1033 : AO4 port map( A => n2558, B => n416, C => n375, D => n2368, Z => 
                           n5139);
   U1034 : AO4 port map( A => n2559, B => n417, C => n2446, D => n2367, Z => 
                           n5140);
   U1035 : AO4 port map( A => n2572, B => n418, C => n2446, D => n2366, Z => 
                           n5141);
   U1037 : AO4 port map( A => n2573, B => n423, C => n375, D => n2365, Z => 
                           n5142);
   U1038 : AO4 port map( A => n2570, B => n424, C => n2446, D => n2364, Z => 
                           n5143);
   U1039 : AO4 port map( A => n2571, B => n425, C => n2446, D => n2363, Z => 
                           n5144);
   U1040 : AO4 port map( A => n2568, B => n426, C => n375, D => n2362, Z => 
                           n5145);
   U1041 : AO4 port map( A => n2569, B => n427, C => n2446, D => n2361, Z => 
                           n5146);
   U1042 : AO4 port map( A => n2566, B => n428, C => n2446, D => n2360, Z => 
                           n5147);
   U1043 : AO4 port map( A => n2567, B => n429, C => n375, D => n2359, Z => 
                           n5148);
   U1044 : AO4 port map( A => n2516, B => n751, C => n2446, D => n2358, Z => 
                           n5149);
   U1045 : AO4 port map( A => n2517, B => n795, C => n2446, D => n2357, Z => 
                           n5150);
   U1046 : AO4 port map( A => n2514, B => n839, C => n375, D => n2356, Z => 
                           n5151);
   U1047 : AO4 port map( A => n2515, B => n883, C => n2446, D => n2355, Z => 
                           n5152);
   U1048 : AO4 port map( A => n2512, B => n430, C => n375, D => n2354, Z => 
                           n5153);
   U1049 : AO4 port map( A => n2513, B => n435, C => n375, D => n2353, Z => 
                           n5154);
   U1050 : AO4 port map( A => n2510, B => n436, C => n375, D => n2352, Z => 
                           n5155);
   U1051 : AO4 port map( A => n2511, B => n437, C => n375, D => n2351, Z => 
                           n5156);
   U1052 : AO4 port map( A => n2524, B => n927, C => n375, D => n2350, Z => 
                           n5157);
   U1053 : AO4 port map( A => n2525, B => n971, C => n375, D => n2349, Z => 
                           n5158);
   U1054 : AO4 port map( A => n2522, B => n1015, C => n375, D => n2348, Z => 
                           n5159);
   U1055 : AO4 port map( A => n2523, B => n1059, C => n375, D => n2347, Z => 
                           n5160);
   U1056 : AO4 port map( A => n2520, B => n438, C => n375, D => n2346, Z => 
                           n5161);
   U1057 : AO4 port map( A => n2521, B => n439, C => n375, D => n2345, Z => 
                           n5162);
   U1058 : AO4 port map( A => n2518, B => n440, C => n375, D => n2344, Z => 
                           n5163);
   U1059 : AO4 port map( A => n2519, B => n441, C => n375, D => n2343, Z => 
                           n5164);
   U1060 : AO4 port map( A => n2532, B => n1103, C => n375, D => n2342, Z => 
                           n5165);
   U1061 : AO4 port map( A => n2533, B => n1147, C => n375, D => n2341, Z => 
                           n5166);
   U1062 : AO4 port map( A => n2530, B => n1191, C => n375, D => n2340, Z => 
                           n5167);
   U1063 : AO4 port map( A => n2531, B => n1235, C => n375, D => n2339, Z => 
                           n5168);
   U1064 : AO4 port map( A => n2528, B => n442, C => n375, D => n2338, Z => 
                           n5169);
   U1065 : AO4 port map( A => n2529, B => n443, C => n375, D => n2337, Z => 
                           n5170);
   U1066 : AO4 port map( A => n2526, B => n487, C => n375, D => n2336, Z => 
                           n5171);
   U1067 : AO4 port map( A => n2527, B => n531, C => n2446, D => n2335, Z => 
                           n5172);
   U1068 : AO4 port map( A => n2540, B => n1279, C => n2446, D => n2334, Z => 
                           n5173);
   U1069 : AO4 port map( A => n2541, B => n1323, C => n2446, D => n2333, Z => 
                           n5174);
   U1070 : AO4 port map( A => n2538, B => n1367, C => n2446, D => n2332, Z => 
                           n5175);
   U1071 : AO4 port map( A => n2539, B => n1411, C => n2446, D => n2331, Z => 
                           n5176);
   U1072 : AO4 port map( A => n2536, B => n575, C => n2446, D => n2330, Z => 
                           n5177);
   U1073 : AO4 port map( A => n2537, B => n619, C => n2446, D => n2329, Z => 
                           n5178);
   U1074 : AO4 port map( A => n2534, B => n663, C => n2446, D => n2328, Z => 
                           n5179);
   U1075 : AO4 port map( A => n2535, B => n707, C => n2446, D => n2327, Z => 
                           n5180);
   U1076 : AO4 port map( A => n2620, B => n390, C => n374, D => n2382, Z => 
                           n5637);
   U1077 : AO4 port map( A => n2621, B => n399, C => n374, D => n2381, Z => 
                           n5638);
   U1078 : AO4 port map( A => n2618, B => n400, C => n374, D => n2380, Z => 
                           n5639);
   U1079 : AO4 port map( A => n2619, B => n401, C => n2454, D => n2379, Z => 
                           n5640);
   U1081 : AO4 port map( A => n2616, B => n402, C => n2454, D => n2378, Z => 
                           n5641);
   U1082 : AO4 port map( A => n2617, B => n403, C => n2454, D => n2377, Z => 
                           n5642);
   U1083 : AO4 port map( A => n2614, B => n404, C => n2454, D => n2376, Z => 
                           n5643);
   U1084 : AO4 port map( A => n2615, B => n405, C => n2454, D => n2375, Z => 
                           n5644);
   U1085 : AO4 port map( A => n2628, B => n406, C => n2454, D => n2374, Z => 
                           n5645);
   U1086 : AO4 port map( A => n2629, B => n411, C => n2454, D => n2373, Z => 
                           n5646);
   U1087 : AO4 port map( A => n2626, B => n412, C => n2454, D => n2372, Z => 
                           n5647);
   U1088 : AO4 port map( A => n2627, B => n413, C => n2454, D => n2371, Z => 
                           n5648);
   U1089 : AO4 port map( A => n2624, B => n414, C => n2454, D => n2370, Z => 
                           n5649);
   U1090 : AO4 port map( A => n2625, B => n415, C => n2454, D => n2369, Z => 
                           n5650);
   U1091 : AO4 port map( A => n2622, B => n416, C => n374, D => n2368, Z => 
                           n5651);
   U1092 : AO4 port map( A => n2623, B => n417, C => n2454, D => n2367, Z => 
                           n5652);
   U1093 : AO4 port map( A => n2636, B => n418, C => n374, D => n2366, Z => 
                           n5653);
   U1094 : AO4 port map( A => n2637, B => n423, C => n2454, D => n2365, Z => 
                           n5654);
   U1095 : AO4 port map( A => n2634, B => n424, C => n374, D => n2364, Z => 
                           n5655);
   U1096 : AO4 port map( A => n2635, B => n425, C => n2454, D => n2363, Z => 
                           n5656);
   U1097 : AO4 port map( A => n2632, B => n426, C => n374, D => n2362, Z => 
                           n5657);
   U1098 : AO4 port map( A => n2633, B => n427, C => n2454, D => n2361, Z => 
                           n5658);
   U1099 : AO4 port map( A => n2630, B => n428, C => n2454, D => n2360, Z => 
                           n5659);
   U1100 : AO4 port map( A => n2631, B => n429, C => n2454, D => n2359, Z => 
                           n5660);
   U1101 : AO4 port map( A => n2580, B => n751, C => n2454, D => n2358, Z => 
                           n5661);
   U1102 : AO4 port map( A => n2581, B => n795, C => n2454, D => n2357, Z => 
                           n5662);
   U1103 : AO4 port map( A => n2578, B => n839, C => n2454, D => n2356, Z => 
                           n5663);
   U1104 : AO4 port map( A => n2579, B => n883, C => n2454, D => n2355, Z => 
                           n5664);
   U1105 : AO4 port map( A => n2576, B => n430, C => n374, D => n2354, Z => 
                           n5665);
   U1106 : AO4 port map( A => n2577, B => n435, C => n2454, D => n2353, Z => 
                           n5666);
   U1107 : AO4 port map( A => n2574, B => n436, C => n2454, D => n2352, Z => 
                           n5667);
   U1108 : AO4 port map( A => n2575, B => n437, C => n374, D => n2351, Z => 
                           n5668);
   U1109 : AO4 port map( A => n2588, B => n927, C => n2454, D => n2350, Z => 
                           n5669);
   U1110 : AO4 port map( A => n2589, B => n971, C => n2454, D => n2349, Z => 
                           n5670);
   U1111 : AO4 port map( A => n2586, B => n1015, C => n374, D => n2348, Z => 
                           n5671);
   U1112 : AO4 port map( A => n2587, B => n1059, C => n374, D => n2347, Z => 
                           n5672);
   U1113 : AO4 port map( A => n2584, B => n438, C => n374, D => n2346, Z => 
                           n5673);
   U1114 : AO4 port map( A => n2585, B => n439, C => n374, D => n2345, Z => 
                           n5674);
   U1115 : AO4 port map( A => n2582, B => n440, C => n374, D => n2344, Z => 
                           n5675);
   U1116 : AO4 port map( A => n2583, B => n441, C => n374, D => n2343, Z => 
                           n5676);
   U1117 : AO4 port map( A => n2596, B => n1103, C => n2454, D => n2342, Z => 
                           n5677);
   U1118 : AO4 port map( A => n2597, B => n1147, C => n2454, D => n2341, Z => 
                           n5678);
   U1119 : AO4 port map( A => n2594, B => n1191, C => n374, D => n2340, Z => 
                           n5679);
   U1120 : AO4 port map( A => n2595, B => n1235, C => n374, D => n2339, Z => 
                           n5680);
   U1121 : AO4 port map( A => n2592, B => n442, C => n374, D => n2338, Z => 
                           n5681);
   U1122 : AO4 port map( A => n2593, B => n443, C => n374, D => n2337, Z => 
                           n5682);
   U1123 : AO4 port map( A => n2590, B => n487, C => n374, D => n2336, Z => 
                           n5683);
   U1125 : AO4 port map( A => n2591, B => n531, C => n374, D => n2335, Z => 
                           n5684);
   U1126 : AO4 port map( A => n2604, B => n1279, C => n374, D => n2334, Z => 
                           n5685);
   U1127 : AO4 port map( A => n2605, B => n1323, C => n374, D => n2333, Z => 
                           n5686);
   U1128 : AO4 port map( A => n2602, B => n1367, C => n374, D => n2332, Z => 
                           n5687);
   U1129 : AO4 port map( A => n2603, B => n1411, C => n374, D => n2331, Z => 
                           n5688);
   U1130 : AO4 port map( A => n2600, B => n575, C => n374, D => n2330, Z => 
                           n5689);
   U1131 : AO4 port map( A => n2601, B => n619, C => n374, D => n2329, Z => 
                           n5690);
   U1132 : AO4 port map( A => n2598, B => n663, C => n374, D => n2328, Z => 
                           n5691);
   U1133 : AO4 port map( A => n2599, B => n707, C => n374, D => n2327, Z => 
                           n5692);
   U1134 : AO4 port map( A => n2684, B => n390, C => n351, D => n2382, Z => 
                           n6149);
   U1135 : AO4 port map( A => n2685, B => n399, C => n351, D => n2381, Z => 
                           n6150);
   U1136 : AO4 port map( A => n2682, B => n400, C => n351, D => n2380, Z => 
                           n6151);
   U1137 : AO4 port map( A => n2683, B => n401, C => n2462, D => n2379, Z => 
                           n6152);
   U1138 : AO4 port map( A => n2680, B => n402, C => n2462, D => n2378, Z => 
                           n6153);
   U1139 : AO4 port map( A => n2681, B => n403, C => n2462, D => n2377, Z => 
                           n6154);
   U1140 : AO4 port map( A => n2678, B => n404, C => n2462, D => n2376, Z => 
                           n6155);
   U1141 : AO4 port map( A => n2679, B => n405, C => n2462, D => n2375, Z => 
                           n6156);
   U1142 : AO4 port map( A => n2692, B => n406, C => n2462, D => n2374, Z => 
                           n6157);
   U1143 : AO4 port map( A => n2693, B => n411, C => n2462, D => n2373, Z => 
                           n6158);
   U1144 : AO4 port map( A => n2690, B => n412, C => n2462, D => n2372, Z => 
                           n6159);
   U1145 : AO4 port map( A => n2691, B => n413, C => n2462, D => n2371, Z => 
                           n6160);
   U1146 : AO4 port map( A => n2688, B => n414, C => n2462, D => n2370, Z => 
                           n6161);
   U1147 : AO4 port map( A => n2689, B => n415, C => n2462, D => n2369, Z => 
                           n6162);
   U1148 : AO4 port map( A => n2686, B => n416, C => n351, D => n2368, Z => 
                           n6163);
   U1149 : AO4 port map( A => n2687, B => n417, C => n2462, D => n2367, Z => 
                           n6164);
   U1150 : AO4 port map( A => n2700, B => n418, C => n351, D => n2366, Z => 
                           n6165);
   U1151 : AO4 port map( A => n2701, B => n423, C => n2462, D => n2365, Z => 
                           n6166);
   U1152 : AO4 port map( A => n2698, B => n424, C => n351, D => n2364, Z => 
                           n6167);
   U1153 : AO4 port map( A => n2699, B => n425, C => n2462, D => n2363, Z => 
                           n6168);
   U1154 : AO4 port map( A => n2696, B => n426, C => n351, D => n2362, Z => 
                           n6169);
   U1155 : AO4 port map( A => n2697, B => n427, C => n2462, D => n2361, Z => 
                           n6170);
   U1156 : AO4 port map( A => n2694, B => n428, C => n2462, D => n2360, Z => 
                           n6171);
   U1157 : AO4 port map( A => n2695, B => n429, C => n2462, D => n2359, Z => 
                           n6172);
   U1158 : AO4 port map( A => n2644, B => n751, C => n2462, D => n2358, Z => 
                           n6173);
   U1159 : AO4 port map( A => n2645, B => n795, C => n2462, D => n2357, Z => 
                           n6174);
   U1160 : AO4 port map( A => n2642, B => n839, C => n2462, D => n2356, Z => 
                           n6175);
   U1161 : AO4 port map( A => n2643, B => n883, C => n2462, D => n2355, Z => 
                           n6176);
   U1162 : AO4 port map( A => n2640, B => n430, C => n351, D => n2354, Z => 
                           n6177);
   U1163 : AO4 port map( A => n2641, B => n435, C => n2462, D => n2353, Z => 
                           n6178);
   U1164 : AO4 port map( A => n2638, B => n436, C => n2462, D => n2352, Z => 
                           n6179);
   U1165 : AO4 port map( A => n2639, B => n437, C => n351, D => n2351, Z => 
                           n6180);
   U1166 : AO4 port map( A => n2652, B => n927, C => n2462, D => n2350, Z => 
                           n6181);
   U1167 : AO4 port map( A => n2653, B => n971, C => n2462, D => n2349, Z => 
                           n6182);
   U1169 : AO4 port map( A => n2650, B => n1015, C => n351, D => n2348, Z => 
                           n6183);
   U1170 : AO4 port map( A => n2651, B => n1059, C => n351, D => n2347, Z => 
                           n6184);
   U1171 : AO4 port map( A => n2648, B => n438, C => n351, D => n2346, Z => 
                           n6185);
   U1172 : AO4 port map( A => n2649, B => n439, C => n351, D => n2345, Z => 
                           n6186);
   U1173 : AO4 port map( A => n2646, B => n440, C => n351, D => n2344, Z => 
                           n6187);
   U1174 : AO4 port map( A => n2647, B => n441, C => n351, D => n2343, Z => 
                           n6188);
   U1175 : AO4 port map( A => n2660, B => n1103, C => n2462, D => n2342, Z => 
                           n6189);
   U1176 : AO4 port map( A => n2661, B => n1147, C => n2462, D => n2341, Z => 
                           n6190);
   U1177 : AO4 port map( A => n2658, B => n1191, C => n351, D => n2340, Z => 
                           n6191);
   U1178 : AO4 port map( A => n2659, B => n1235, C => n351, D => n2339, Z => 
                           n6192);
   U1179 : AO4 port map( A => n2656, B => n442, C => n351, D => n2338, Z => 
                           n6193);
   U1180 : AO4 port map( A => n2657, B => n443, C => n351, D => n2337, Z => 
                           n6194);
   U1181 : AO4 port map( A => n2654, B => n487, C => n351, D => n2336, Z => 
                           n6195);
   U1182 : AO4 port map( A => n2655, B => n531, C => n351, D => n2335, Z => 
                           n6196);
   U1183 : AO4 port map( A => n2668, B => n1279, C => n351, D => n2334, Z => 
                           n6197);
   U1184 : AO4 port map( A => n2669, B => n1323, C => n351, D => n2333, Z => 
                           n6198);
   U1185 : AO4 port map( A => n2666, B => n1367, C => n351, D => n2332, Z => 
                           n6199);
   U1186 : AO4 port map( A => n2667, B => n1411, C => n351, D => n2331, Z => 
                           n6200);
   U1187 : AO4 port map( A => n2664, B => n575, C => n351, D => n2330, Z => 
                           n6201);
   U1188 : AO4 port map( A => n2665, B => n619, C => n351, D => n2329, Z => 
                           n6202);
   U1189 : AO4 port map( A => n2662, B => n663, C => n351, D => n2328, Z => 
                           n6203);
   U1190 : AO4 port map( A => n2663, B => n707, C => n351, D => n2327, Z => 
                           n6204);
   U1191 : AO4 port map( A => n2740, B => n378, C => n2309, D => n2390, Z => 
                           n4605);
   U1192 : AO4 port map( A => n2741, B => n383, C => n2309, D => n2389, Z => 
                           n4606);
   U1193 : AO4 port map( A => n2738, B => n384, C => n2309, D => n2388, Z => 
                           n4607);
   U1194 : AO4 port map( A => n2739, B => n385, C => n2309, D => n2387, Z => 
                           n4608);
   U1195 : AO4 port map( A => n2736, B => n386, C => n2309, D => n2386, Z => 
                           n4609);
   U1196 : AO4 port map( A => n2737, B => n387, C => n2309, D => n2385, Z => 
                           n4610);
   U1197 : AO4 port map( A => n2734, B => n388, C => n2309, D => n2384, Z => 
                           n4611);
   U1198 : AO4 port map( A => n2735, B => n389, C => n2309, D => n2383, Z => 
                           n4612);
   U1199 : AO4 port map( A => n2748, B => n390, C => n2309, D => n2382, Z => 
                           n4613);
   U1200 : AO4 port map( A => n2749, B => n399, C => n2309, D => n2381, Z => 
                           n4614);
   U1201 : AO4 port map( A => n2746, B => n400, C => n2309, D => n2380, Z => 
                           n4615);
   U1202 : AO4 port map( A => n2747, B => n401, C => n2309, D => n2379, Z => 
                           n4616);
   U1203 : AO4 port map( A => n2744, B => n402, C => n2309, D => n2378, Z => 
                           n4617);
   U1204 : AO4 port map( A => n2745, B => n403, C => n2309, D => n2377, Z => 
                           n4618);
   U1205 : AO4 port map( A => n2742, B => n404, C => n2309, D => n2376, Z => 
                           n4619);
   U1206 : AO4 port map( A => n2743, B => n405, C => n2309, D => n2375, Z => 
                           n4620);
   U1207 : AO4 port map( A => n2756, B => n406, C => n353, D => n2374, Z => 
                           n4621);
   U1208 : AO4 port map( A => n2757, B => n411, C => n2309, D => n2373, Z => 
                           n4622);
   U1209 : AO4 port map( A => n2754, B => n412, C => n2309, D => n2372, Z => 
                           n4623);
   U1210 : AO4 port map( A => n2755, B => n413, C => n2309, D => n2371, Z => 
                           n4624);
   U1211 : AO4 port map( A => n2752, B => n414, C => n353, D => n2370, Z => 
                           n4625);
   U1213 : AO4 port map( A => n2753, B => n415, C => n2309, D => n2369, Z => 
                           n4626);
   U1214 : AO4 port map( A => n2750, B => n416, C => n353, D => n2368, Z => 
                           n4627);
   U1215 : AO4 port map( A => n2751, B => n417, C => n353, D => n2367, Z => 
                           n4628);
   U1216 : AO4 port map( A => n2764, B => n418, C => n353, D => n2366, Z => 
                           n4629);
   U1217 : AO4 port map( A => n2765, B => n423, C => n353, D => n2365, Z => 
                           n4630);
   U1218 : AO4 port map( A => n2762, B => n424, C => n353, D => n2364, Z => 
                           n4631);
   U1219 : AO4 port map( A => n2763, B => n425, C => n353, D => n2363, Z => 
                           n4632);
   U1220 : AO4 port map( A => n2760, B => n426, C => n353, D => n2362, Z => 
                           n4633);
   U1221 : AO4 port map( A => n2761, B => n427, C => n353, D => n2361, Z => 
                           n4634);
   U1222 : AO4 port map( A => n2758, B => n428, C => n353, D => n2360, Z => 
                           n4635);
   U1223 : AO4 port map( A => n2759, B => n429, C => n353, D => n2359, Z => 
                           n4636);
   U1224 : AO4 port map( A => n2708, B => n751, C => n353, D => n2358, Z => 
                           n4637);
   U1225 : AO4 port map( A => n2709, B => n795, C => n353, D => n2357, Z => 
                           n4638);
   U1226 : AO4 port map( A => n2706, B => n839, C => n353, D => n2356, Z => 
                           n4639);
   U1227 : AO4 port map( A => n2707, B => n883, C => n353, D => n2355, Z => 
                           n4640);
   U1228 : AO4 port map( A => n2704, B => n430, C => n353, D => n2354, Z => 
                           n4641);
   U1229 : AO4 port map( A => n2705, B => n435, C => n353, D => n2353, Z => 
                           n4642);
   U1230 : AO4 port map( A => n2702, B => n436, C => n353, D => n2352, Z => 
                           n4643);
   U1231 : AO4 port map( A => n2703, B => n437, C => n353, D => n2351, Z => 
                           n4644);
   U1232 : AO4 port map( A => n2716, B => n927, C => n353, D => n2350, Z => 
                           n4645);
   U1233 : AO4 port map( A => n2717, B => n971, C => n353, D => n2349, Z => 
                           n4646);
   U1234 : AO4 port map( A => n2714, B => n1015, C => n353, D => n2348, Z => 
                           n4647);
   U1235 : AO4 port map( A => n2715, B => n1059, C => n353, D => n2347, Z => 
                           n4648);
   U1236 : AO4 port map( A => n2712, B => n438, C => n353, D => n2346, Z => 
                           n4649);
   U1237 : AO4 port map( A => n2713, B => n439, C => n353, D => n2345, Z => 
                           n4650);
   U1238 : AO4 port map( A => n2710, B => n440, C => n2309, D => n2344, Z => 
                           n4651);
   U1239 : AO4 port map( A => n2711, B => n441, C => n2309, D => n2343, Z => 
                           n4652);
   U1240 : AO4 port map( A => n2724, B => n1103, C => n2309, D => n2342, Z => 
                           n4653);
   U1241 : AO4 port map( A => n2725, B => n1147, C => n2309, D => n2341, Z => 
                           n4654);
   U1242 : AO4 port map( A => n2722, B => n1191, C => n2309, D => n2340, Z => 
                           n4655);
   U1243 : AO4 port map( A => n2723, B => n1235, C => n353, D => n2339, Z => 
                           n4656);
   U1244 : AO4 port map( A => n2720, B => n442, C => n2309, D => n2338, Z => 
                           n4657);
   U1245 : AO4 port map( A => n2721, B => n443, C => n2309, D => n2337, Z => 
                           n4658);
   U1246 : AO4 port map( A => n2718, B => n487, C => n353, D => n2336, Z => 
                           n4659);
   U1247 : AO4 port map( A => n2719, B => n531, C => n2309, D => n2335, Z => 
                           n4660);
   U1248 : AO4 port map( A => n2732, B => n1279, C => n2309, D => n2334, Z => 
                           n4661);
   U1249 : AO4 port map( A => n2733, B => n1323, C => n353, D => n2333, Z => 
                           n4662);
   U1250 : AO4 port map( A => n2730, B => n1367, C => n2309, D => n2332, Z => 
                           n4663);
   U1251 : AO4 port map( A => n2731, B => n1411, C => n2309, D => n2331, Z => 
                           n4664);
   U1252 : AO4 port map( A => n2728, B => n575, C => n353, D => n2330, Z => 
                           n4665);
   U1253 : AO4 port map( A => n2729, B => n619, C => n2309, D => n2329, Z => 
                           n4666);
   U1254 : AO4 port map( A => n2726, B => n663, C => n2309, D => n2328, Z => 
                           n4667);
   U1255 : AO4 port map( A => n2727, B => n707, C => n353, D => n2327, Z => 
                           n4668);
   U1257 : AO4 port map( A => n2812, B => n390, C => n373, D => n2382, Z => 
                           n5189);
   U1258 : AO4 port map( A => n2813, B => n399, C => n2447, D => n2381, Z => 
                           n5190);
   U1259 : AO4 port map( A => n2810, B => n400, C => n373, D => n2380, Z => 
                           n5191);
   U1260 : AO4 port map( A => n2811, B => n401, C => n2447, D => n2379, Z => 
                           n5192);
   U1261 : AO4 port map( A => n2808, B => n402, C => n373, D => n2378, Z => 
                           n5193);
   U1262 : AO4 port map( A => n2809, B => n403, C => n2447, D => n2377, Z => 
                           n5194);
   U1263 : AO4 port map( A => n2806, B => n404, C => n373, D => n2376, Z => 
                           n5195);
   U1264 : AO4 port map( A => n2807, B => n405, C => n2447, D => n2375, Z => 
                           n5196);
   U1265 : AO4 port map( A => n2820, B => n406, C => n373, D => n2374, Z => 
                           n5197);
   U1266 : AO4 port map( A => n2821, B => n411, C => n2447, D => n2373, Z => 
                           n5198);
   U1267 : AO4 port map( A => n2818, B => n412, C => n2447, D => n2372, Z => 
                           n5199);
   U1268 : AO4 port map( A => n2819, B => n413, C => n2447, D => n2371, Z => 
                           n5200);
   U1269 : AO4 port map( A => n2816, B => n414, C => n2447, D => n2370, Z => 
                           n5201);
   U1270 : AO4 port map( A => n2817, B => n415, C => n2447, D => n2369, Z => 
                           n5202);
   U1271 : AO4 port map( A => n2814, B => n416, C => n373, D => n2368, Z => 
                           n5203);
   U1272 : AO4 port map( A => n2815, B => n417, C => n2447, D => n2367, Z => 
                           n5204);
   U1273 : AO4 port map( A => n2828, B => n418, C => n2447, D => n2366, Z => 
                           n5205);
   U1274 : AO4 port map( A => n2829, B => n423, C => n373, D => n2365, Z => 
                           n5206);
   U1275 : AO4 port map( A => n2826, B => n424, C => n2447, D => n2364, Z => 
                           n5207);
   U1276 : AO4 port map( A => n2827, B => n425, C => n2447, D => n2363, Z => 
                           n5208);
   U1277 : AO4 port map( A => n2824, B => n426, C => n373, D => n2362, Z => 
                           n5209);
   U1278 : AO4 port map( A => n2825, B => n427, C => n2447, D => n2361, Z => 
                           n5210);
   U1279 : AO4 port map( A => n2822, B => n428, C => n2447, D => n2360, Z => 
                           n5211);
   U1280 : AO4 port map( A => n2823, B => n429, C => n373, D => n2359, Z => 
                           n5212);
   U1281 : AO4 port map( A => n2772, B => n751, C => n2447, D => n2358, Z => 
                           n5213);
   U1282 : AO4 port map( A => n2773, B => n795, C => n2447, D => n2357, Z => 
                           n5214);
   U1283 : AO4 port map( A => n2770, B => n839, C => n373, D => n2356, Z => 
                           n5215);
   U1284 : AO4 port map( A => n2771, B => n883, C => n2447, D => n2355, Z => 
                           n5216);
   U1285 : AO4 port map( A => n2768, B => n430, C => n373, D => n2354, Z => 
                           n5217);
   U1286 : AO4 port map( A => n2769, B => n435, C => n373, D => n2353, Z => 
                           n5218);
   U1287 : AO4 port map( A => n2766, B => n436, C => n373, D => n2352, Z => 
                           n5219);
   U1288 : AO4 port map( A => n2767, B => n437, C => n373, D => n2351, Z => 
                           n5220);
   U1289 : AO4 port map( A => n2780, B => n927, C => n373, D => n2350, Z => 
                           n5221);
   U1290 : AO4 port map( A => n2781, B => n971, C => n373, D => n2349, Z => 
                           n5222);
   U1291 : AO4 port map( A => n2778, B => n1015, C => n373, D => n2348, Z => 
                           n5223);
   U1292 : AO4 port map( A => n2779, B => n1059, C => n373, D => n2347, Z => 
                           n5224);
   U1293 : AO4 port map( A => n2776, B => n438, C => n373, D => n2346, Z => 
                           n5225);
   U1294 : AO4 port map( A => n2777, B => n439, C => n373, D => n2345, Z => 
                           n5226);
   U1295 : AO4 port map( A => n2774, B => n440, C => n373, D => n2344, Z => 
                           n5227);
   U1296 : AO4 port map( A => n2775, B => n441, C => n373, D => n2343, Z => 
                           n5228);
   U1297 : AO4 port map( A => n2788, B => n1103, C => n373, D => n2342, Z => 
                           n5229);
   U1298 : AO4 port map( A => n2789, B => n1147, C => n373, D => n2341, Z => 
                           n5230);
   U1299 : AO4 port map( A => n2786, B => n1191, C => n373, D => n2340, Z => 
                           n5231);
   U1301 : AO4 port map( A => n2787, B => n1235, C => n373, D => n2339, Z => 
                           n5232);
   U1302 : AO4 port map( A => n2784, B => n442, C => n373, D => n2338, Z => 
                           n5233);
   U1303 : AO4 port map( A => n2785, B => n443, C => n373, D => n2337, Z => 
                           n5234);
   U1304 : AO4 port map( A => n2782, B => n487, C => n373, D => n2336, Z => 
                           n5235);
   U1305 : AO4 port map( A => n2783, B => n531, C => n2447, D => n2335, Z => 
                           n5236);
   U1306 : AO4 port map( A => n2796, B => n1279, C => n2447, D => n2334, Z => 
                           n5237);
   U1307 : AO4 port map( A => n2797, B => n1323, C => n2447, D => n2333, Z => 
                           n5238);
   U1308 : AO4 port map( A => n2794, B => n1367, C => n2447, D => n2332, Z => 
                           n5239);
   U1309 : AO4 port map( A => n2795, B => n1411, C => n2447, D => n2331, Z => 
                           n5240);
   U1310 : AO4 port map( A => n2792, B => n575, C => n2447, D => n2330, Z => 
                           n5241);
   U1311 : AO4 port map( A => n2793, B => n619, C => n2447, D => n2329, Z => 
                           n5242);
   U1312 : AO4 port map( A => n2790, B => n663, C => n2447, D => n2328, Z => 
                           n5243);
   U1313 : AO4 port map( A => n2791, B => n707, C => n2447, D => n2327, Z => 
                           n5244);
   U1314 : AO4 port map( A => n2876, B => n390, C => n372, D => n2382, Z => 
                           n5701);
   U1315 : AO4 port map( A => n2877, B => n399, C => n2455, D => n2381, Z => 
                           n5702);
   U1316 : AO4 port map( A => n2874, B => n400, C => n372, D => n2380, Z => 
                           n5703);
   U1317 : AO4 port map( A => n2875, B => n401, C => n2455, D => n2379, Z => 
                           n5704);
   U1318 : AO4 port map( A => n2872, B => n402, C => n372, D => n2378, Z => 
                           n5705);
   U1319 : AO4 port map( A => n2873, B => n403, C => n2455, D => n2377, Z => 
                           n5706);
   U1320 : AO4 port map( A => n2870, B => n404, C => n372, D => n2376, Z => 
                           n5707);
   U1321 : AO4 port map( A => n2871, B => n405, C => n2455, D => n2375, Z => 
                           n5708);
   U1322 : AO4 port map( A => n2884, B => n406, C => n372, D => n2374, Z => 
                           n5709);
   U1323 : AO4 port map( A => n2885, B => n411, C => n2455, D => n2373, Z => 
                           n5710);
   U1324 : AO4 port map( A => n2882, B => n412, C => n2455, D => n2372, Z => 
                           n5711);
   U1325 : AO4 port map( A => n2883, B => n413, C => n2455, D => n2371, Z => 
                           n5712);
   U1326 : AO4 port map( A => n2880, B => n414, C => n2455, D => n2370, Z => 
                           n5713);
   U1327 : AO4 port map( A => n2881, B => n415, C => n2455, D => n2369, Z => 
                           n5714);
   U1328 : AO4 port map( A => n2878, B => n416, C => n372, D => n2368, Z => 
                           n5715);
   U1329 : AO4 port map( A => n2879, B => n417, C => n2455, D => n2367, Z => 
                           n5716);
   U1330 : AO4 port map( A => n2892, B => n418, C => n2455, D => n2366, Z => 
                           n5717);
   U1331 : AO4 port map( A => n2893, B => n423, C => n372, D => n2365, Z => 
                           n5718);
   U1332 : AO4 port map( A => n2890, B => n424, C => n2455, D => n2364, Z => 
                           n5719);
   U1333 : AO4 port map( A => n2891, B => n425, C => n2455, D => n2363, Z => 
                           n5720);
   U1334 : AO4 port map( A => n2888, B => n426, C => n372, D => n2362, Z => 
                           n5721);
   U1335 : AO4 port map( A => n2889, B => n427, C => n2455, D => n2361, Z => 
                           n5722);
   U1336 : AO4 port map( A => n2886, B => n428, C => n2455, D => n2360, Z => 
                           n5723);
   U1337 : AO4 port map( A => n2887, B => n429, C => n372, D => n2359, Z => 
                           n5724);
   U1338 : AO4 port map( A => n2836, B => n751, C => n2455, D => n2358, Z => 
                           n5725);
   U1339 : AO4 port map( A => n2837, B => n795, C => n2455, D => n2357, Z => 
                           n5726);
   U1340 : AO4 port map( A => n2834, B => n839, C => n372, D => n2356, Z => 
                           n5727);
   U1341 : AO4 port map( A => n2835, B => n883, C => n2455, D => n2355, Z => 
                           n5728);
   U1342 : AO4 port map( A => n2832, B => n430, C => n372, D => n2354, Z => 
                           n5729);
   U1343 : AO4 port map( A => n2833, B => n435, C => n372, D => n2353, Z => 
                           n5730);
   U1345 : AO4 port map( A => n2830, B => n436, C => n372, D => n2352, Z => 
                           n5731);
   U1346 : AO4 port map( A => n2831, B => n437, C => n372, D => n2351, Z => 
                           n5732);
   U1347 : AO4 port map( A => n2844, B => n927, C => n372, D => n2350, Z => 
                           n5733);
   U1348 : AO4 port map( A => n2845, B => n971, C => n372, D => n2349, Z => 
                           n5734);
   U1349 : AO4 port map( A => n2842, B => n1015, C => n372, D => n2348, Z => 
                           n5735);
   U1350 : AO4 port map( A => n2843, B => n1059, C => n372, D => n2347, Z => 
                           n5736);
   U1351 : AO4 port map( A => n2840, B => n438, C => n372, D => n2346, Z => 
                           n5737);
   U1352 : AO4 port map( A => n2841, B => n439, C => n372, D => n2345, Z => 
                           n5738);
   U1353 : AO4 port map( A => n2838, B => n440, C => n372, D => n2344, Z => 
                           n5739);
   U1354 : AO4 port map( A => n2839, B => n441, C => n372, D => n2343, Z => 
                           n5740);
   U1355 : AO4 port map( A => n2852, B => n1103, C => n372, D => n2342, Z => 
                           n5741);
   U1356 : AO4 port map( A => n2853, B => n1147, C => n372, D => n2341, Z => 
                           n5742);
   U1357 : AO4 port map( A => n2850, B => n1191, C => n372, D => n2340, Z => 
                           n5743);
   U1358 : AO4 port map( A => n2851, B => n1235, C => n372, D => n2339, Z => 
                           n5744);
   U1359 : AO4 port map( A => n2848, B => n442, C => n372, D => n2338, Z => 
                           n5745);
   U1360 : AO4 port map( A => n2849, B => n443, C => n372, D => n2337, Z => 
                           n5746);
   U1361 : AO4 port map( A => n2846, B => n487, C => n372, D => n2336, Z => 
                           n5747);
   U1362 : AO4 port map( A => n2847, B => n531, C => n2455, D => n2335, Z => 
                           n5748);
   U1363 : AO4 port map( A => n2860, B => n1279, C => n2455, D => n2334, Z => 
                           n5749);
   U1364 : AO4 port map( A => n2861, B => n1323, C => n2455, D => n2333, Z => 
                           n5750);
   U1365 : AO4 port map( A => n2858, B => n1367, C => n2455, D => n2332, Z => 
                           n5751);
   U1366 : AO4 port map( A => n2859, B => n1411, C => n2455, D => n2331, Z => 
                           n5752);
   U1367 : AO4 port map( A => n2856, B => n575, C => n2455, D => n2330, Z => 
                           n5753);
   U1368 : AO4 port map( A => n2857, B => n619, C => n2455, D => n2329, Z => 
                           n5754);
   U1369 : AO4 port map( A => n2854, B => n663, C => n2455, D => n2328, Z => 
                           n5755);
   U1370 : AO4 port map( A => n2855, B => n707, C => n2455, D => n2327, Z => 
                           n5756);
   U1371 : AO4 port map( A => n2940, B => n390, C => n350, D => n2382, Z => 
                           n6213);
   U1372 : AO4 port map( A => n2941, B => n399, C => n2463, D => n2381, Z => 
                           n6214);
   U1373 : AO4 port map( A => n2938, B => n400, C => n350, D => n2380, Z => 
                           n6215);
   U1374 : AO4 port map( A => n2939, B => n401, C => n2463, D => n2379, Z => 
                           n6216);
   U1375 : AO4 port map( A => n2936, B => n402, C => n350, D => n2378, Z => 
                           n6217);
   U1376 : AO4 port map( A => n2937, B => n403, C => n2463, D => n2377, Z => 
                           n6218);
   U1377 : AO4 port map( A => n2934, B => n404, C => n350, D => n2376, Z => 
                           n6219);
   U1378 : AO4 port map( A => n2935, B => n405, C => n2463, D => n2375, Z => 
                           n6220);
   U1379 : AO4 port map( A => n2948, B => n406, C => n350, D => n2374, Z => 
                           n6221);
   U1380 : AO4 port map( A => n2949, B => n411, C => n2463, D => n2373, Z => 
                           n6222);
   U1381 : AO4 port map( A => n2946, B => n412, C => n2463, D => n2372, Z => 
                           n6223);
   U1382 : AO4 port map( A => n2947, B => n413, C => n2463, D => n2371, Z => 
                           n6224);
   U1383 : AO4 port map( A => n2944, B => n414, C => n2463, D => n2370, Z => 
                           n6225);
   U1384 : AO4 port map( A => n2945, B => n415, C => n2463, D => n2369, Z => 
                           n6226);
   U1385 : AO4 port map( A => n2942, B => n416, C => n350, D => n2368, Z => 
                           n6227);
   U1386 : AO4 port map( A => n2943, B => n417, C => n2463, D => n2367, Z => 
                           n6228);
   U1387 : AO4 port map( A => n2956, B => n418, C => n2463, D => n2366, Z => 
                           n6229);
   U1389 : AO4 port map( A => n2957, B => n423, C => n350, D => n2365, Z => 
                           n6230);
   U1390 : AO4 port map( A => n2954, B => n424, C => n2463, D => n2364, Z => 
                           n6231);
   U1391 : AO4 port map( A => n2955, B => n425, C => n2463, D => n2363, Z => 
                           n6232);
   U1392 : AO4 port map( A => n2952, B => n426, C => n350, D => n2362, Z => 
                           n6233);
   U1393 : AO4 port map( A => n2953, B => n427, C => n2463, D => n2361, Z => 
                           n6234);
   U1394 : AO4 port map( A => n2950, B => n428, C => n2463, D => n2360, Z => 
                           n6235);
   U1395 : AO4 port map( A => n2951, B => n429, C => n350, D => n2359, Z => 
                           n6236);
   U1396 : AO4 port map( A => n2900, B => n751, C => n2463, D => n2358, Z => 
                           n6237);
   U1397 : AO4 port map( A => n2901, B => n795, C => n2463, D => n2357, Z => 
                           n6238);
   U1398 : AO4 port map( A => n2898, B => n839, C => n350, D => n2356, Z => 
                           n6239);
   U1399 : AO4 port map( A => n2899, B => n883, C => n2463, D => n2355, Z => 
                           n6240);
   U1400 : AO4 port map( A => n2896, B => n430, C => n350, D => n2354, Z => 
                           n6241);
   U1401 : AO4 port map( A => n2897, B => n435, C => n350, D => n2353, Z => 
                           n6242);
   U1402 : AO4 port map( A => n2894, B => n436, C => n350, D => n2352, Z => 
                           n6243);
   U1403 : AO4 port map( A => n2895, B => n437, C => n350, D => n2351, Z => 
                           n6244);
   U1404 : AO4 port map( A => n2908, B => n927, C => n350, D => n2350, Z => 
                           n6245);
   U1405 : AO4 port map( A => n2909, B => n971, C => n350, D => n2349, Z => 
                           n6246);
   U1406 : AO4 port map( A => n2906, B => n1015, C => n350, D => n2348, Z => 
                           n6247);
   U1407 : AO4 port map( A => n2907, B => n1059, C => n350, D => n2347, Z => 
                           n6248);
   U1408 : AO4 port map( A => n2904, B => n438, C => n350, D => n2346, Z => 
                           n6249);
   U1409 : AO4 port map( A => n2905, B => n439, C => n350, D => n2345, Z => 
                           n6250);
   U1410 : AO4 port map( A => n2902, B => n440, C => n350, D => n2344, Z => 
                           n6251);
   U1411 : AO4 port map( A => n2903, B => n441, C => n350, D => n2343, Z => 
                           n6252);
   U1412 : AO4 port map( A => n2916, B => n1103, C => n350, D => n2342, Z => 
                           n6253);
   U1413 : AO4 port map( A => n2917, B => n1147, C => n350, D => n2341, Z => 
                           n6254);
   U1414 : AO4 port map( A => n2914, B => n1191, C => n350, D => n2340, Z => 
                           n6255);
   U1415 : AO4 port map( A => n2915, B => n1235, C => n350, D => n2339, Z => 
                           n6256);
   U1416 : AO4 port map( A => n2912, B => n442, C => n350, D => n2338, Z => 
                           n6257);
   U1417 : AO4 port map( A => n2913, B => n443, C => n350, D => n2337, Z => 
                           n6258);
   U1418 : AO4 port map( A => n2910, B => n487, C => n350, D => n2336, Z => 
                           n6259);
   U1419 : AO4 port map( A => n2911, B => n531, C => n2463, D => n2335, Z => 
                           n6260);
   U1420 : AO4 port map( A => n2924, B => n1279, C => n2463, D => n2334, Z => 
                           n6261);
   U1421 : AO4 port map( A => n2925, B => n1323, C => n2463, D => n2333, Z => 
                           n6262);
   U1422 : AO4 port map( A => n2922, B => n1367, C => n2463, D => n2332, Z => 
                           n6263);
   U1423 : AO4 port map( A => n2923, B => n1411, C => n2463, D => n2331, Z => 
                           n6264);
   U1424 : AO4 port map( A => n2920, B => n575, C => n2463, D => n2330, Z => 
                           n6265);
   U1425 : AO4 port map( A => n2921, B => n619, C => n2463, D => n2329, Z => 
                           n6266);
   U1426 : AO4 port map( A => n2918, B => n663, C => n2463, D => n2328, Z => 
                           n6267);
   U1427 : AO4 port map( A => n2919, B => n707, C => n2463, D => n2327, Z => 
                           n6268);
   U1428 : AO4 port map( A => n2996, B => n378, C => n377, D => n2390, Z => 
                           n4669);
   U1429 : AO4 port map( A => n2997, B => n383, C => n2439, D => n2389, Z => 
                           n4670);
   U1430 : AO4 port map( A => n2994, B => n384, C => n2439, D => n2388, Z => 
                           n4671);
   U1431 : AO4 port map( A => n2995, B => n385, C => n2439, D => n2387, Z => 
                           n4672);
   U1433 : AO4 port map( A => n2992, B => n386, C => n377, D => n2386, Z => 
                           n4673);
   U1434 : AO4 port map( A => n2993, B => n387, C => n2439, D => n2385, Z => 
                           n4674);
   U1435 : AO4 port map( A => n2990, B => n388, C => n2439, D => n2384, Z => 
                           n4675);
   U1436 : AO4 port map( A => n2991, B => n389, C => n2439, D => n2383, Z => 
                           n4676);
   U1437 : AO4 port map( A => n3004, B => n390, C => n377, D => n2382, Z => 
                           n4677);
   U1438 : AO4 port map( A => n3005, B => n399, C => n2439, D => n2381, Z => 
                           n4678);
   U1439 : AO4 port map( A => n3002, B => n400, C => n377, D => n2380, Z => 
                           n4679);
   U1440 : AO4 port map( A => n3003, B => n401, C => n2439, D => n2379, Z => 
                           n4680);
   U1441 : AO4 port map( A => n3000, B => n402, C => n377, D => n2378, Z => 
                           n4681);
   U1442 : AO4 port map( A => n3001, B => n403, C => n2439, D => n2377, Z => 
                           n4682);
   U1443 : AO4 port map( A => n2998, B => n404, C => n377, D => n2376, Z => 
                           n4683);
   U1444 : AO4 port map( A => n2999, B => n405, C => n2439, D => n2375, Z => 
                           n4684);
   U1445 : AO4 port map( A => n3012, B => n406, C => n377, D => n2374, Z => 
                           n4685);
   U1446 : AO4 port map( A => n3013, B => n411, C => n2439, D => n2373, Z => 
                           n4686);
   U1447 : AO4 port map( A => n3010, B => n412, C => n2439, D => n2372, Z => 
                           n4687);
   U1448 : AO4 port map( A => n3011, B => n413, C => n2439, D => n2371, Z => 
                           n4688);
   U1449 : AO4 port map( A => n3008, B => n414, C => n2439, D => n2370, Z => 
                           n4689);
   U1450 : AO4 port map( A => n3009, B => n415, C => n2439, D => n2369, Z => 
                           n4690);
   U1451 : AO4 port map( A => n3006, B => n416, C => n377, D => n2368, Z => 
                           n4691);
   U1452 : AO4 port map( A => n3007, B => n417, C => n2439, D => n2367, Z => 
                           n4692);
   U1453 : AO4 port map( A => n3020, B => n418, C => n2439, D => n2366, Z => 
                           n4693);
   U1454 : AO4 port map( A => n3021, B => n423, C => n377, D => n2365, Z => 
                           n4694);
   U1455 : AO4 port map( A => n3018, B => n424, C => n2439, D => n2364, Z => 
                           n4695);
   U1456 : AO4 port map( A => n3019, B => n425, C => n2439, D => n2363, Z => 
                           n4696);
   U1457 : AO4 port map( A => n3016, B => n426, C => n377, D => n2362, Z => 
                           n4697);
   U1458 : AO4 port map( A => n3017, B => n427, C => n2439, D => n2361, Z => 
                           n4698);
   U1459 : AO4 port map( A => n3014, B => n428, C => n2439, D => n2360, Z => 
                           n4699);
   U1460 : AO4 port map( A => n3015, B => n429, C => n377, D => n2359, Z => 
                           n4700);
   U1461 : AO4 port map( A => n2964, B => n751, C => n2439, D => n2358, Z => 
                           n4701);
   U1462 : AO4 port map( A => n2965, B => n795, C => n2439, D => n2357, Z => 
                           n4702);
   U1463 : AO4 port map( A => n2962, B => n839, C => n377, D => n2356, Z => 
                           n4703);
   U1464 : AO4 port map( A => n2963, B => n883, C => n2439, D => n2355, Z => 
                           n4704);
   U1465 : AO4 port map( A => n2960, B => n430, C => n377, D => n2354, Z => 
                           n4705);
   U1466 : AO4 port map( A => n2961, B => n435, C => n377, D => n2353, Z => 
                           n4706);
   U1467 : AO4 port map( A => n2958, B => n436, C => n377, D => n2352, Z => 
                           n4707);
   U1468 : AO4 port map( A => n2959, B => n437, C => n377, D => n2351, Z => 
                           n4708);
   U1469 : AO4 port map( A => n2972, B => n927, C => n377, D => n2350, Z => 
                           n4709);
   U1470 : AO4 port map( A => n2973, B => n971, C => n377, D => n2349, Z => 
                           n4710);
   U1471 : AO4 port map( A => n2970, B => n1015, C => n377, D => n2348, Z => 
                           n4711);
   U1472 : AO4 port map( A => n2971, B => n1059, C => n377, D => n2347, Z => 
                           n4712);
   U1473 : AO4 port map( A => n2968, B => n438, C => n377, D => n2346, Z => 
                           n4713);
   U1474 : AO4 port map( A => n2969, B => n439, C => n377, D => n2345, Z => 
                           n4714);
   U1475 : AO4 port map( A => n2966, B => n440, C => n377, D => n2344, Z => 
                           n4715);
   U1477 : AO4 port map( A => n2967, B => n441, C => n377, D => n2343, Z => 
                           n4716);
   U1478 : AO4 port map( A => n2980, B => n1103, C => n377, D => n2342, Z => 
                           n4717);
   U1479 : AO4 port map( A => n2981, B => n1147, C => n377, D => n2341, Z => 
                           n4718);
   U1480 : AO4 port map( A => n2978, B => n1191, C => n377, D => n2340, Z => 
                           n4719);
   U1481 : AO4 port map( A => n2979, B => n1235, C => n377, D => n2339, Z => 
                           n4720);
   U1482 : AO4 port map( A => n2976, B => n442, C => n377, D => n2338, Z => 
                           n4721);
   U1483 : AO4 port map( A => n2977, B => n443, C => n377, D => n2337, Z => 
                           n4722);
   U1484 : AO4 port map( A => n2974, B => n487, C => n377, D => n2336, Z => 
                           n4723);
   U1485 : AO4 port map( A => n2975, B => n531, C => n2439, D => n2335, Z => 
                           n4724);
   U1486 : AO4 port map( A => n2988, B => n1279, C => n2439, D => n2334, Z => 
                           n4725);
   U1487 : AO4 port map( A => n2989, B => n1323, C => n2439, D => n2333, Z => 
                           n4726);
   U1488 : AO4 port map( A => n2986, B => n1367, C => n2439, D => n2332, Z => 
                           n4727);
   U1489 : AO4 port map( A => n2987, B => n1411, C => n2439, D => n2331, Z => 
                           n4728);
   U1490 : AO4 port map( A => n2984, B => n575, C => n2439, D => n2330, Z => 
                           n4729);
   U1491 : AO4 port map( A => n2985, B => n619, C => n2439, D => n2329, Z => 
                           n4730);
   U1492 : AO4 port map( A => n2982, B => n663, C => n2439, D => n2328, Z => 
                           n4731);
   U1493 : AO4 port map( A => n2983, B => n707, C => n2439, D => n2327, Z => 
                           n4732);
   U1494 : AO4 port map( A => n3068, B => n390, C => n2448, D => n2382, Z => 
                           n5253);
   U1495 : AO4 port map( A => n3069, B => n399, C => n2448, D => n2381, Z => 
                           n5254);
   U1496 : AO4 port map( A => n3066, B => n400, C => n2448, D => n2380, Z => 
                           n5255);
   U1497 : AO4 port map( A => n3067, B => n401, C => n2448, D => n2379, Z => 
                           n5256);
   U1498 : AO4 port map( A => n3064, B => n402, C => n2448, D => n2378, Z => 
                           n5257);
   U1499 : AO4 port map( A => n3065, B => n403, C => n2448, D => n2377, Z => 
                           n5258);
   U1500 : AO4 port map( A => n3062, B => n404, C => n2448, D => n2376, Z => 
                           n5259);
   U1501 : AO4 port map( A => n3063, B => n405, C => n2448, D => n2375, Z => 
                           n5260);
   U1502 : AO4 port map( A => n3076, B => n406, C => n371, D => n2374, Z => 
                           n5261);
   U1503 : AO4 port map( A => n3077, B => n411, C => n2448, D => n2373, Z => 
                           n5262);
   U1504 : AO4 port map( A => n3074, B => n412, C => n2448, D => n2372, Z => 
                           n5263);
   U1505 : AO4 port map( A => n3075, B => n413, C => n2448, D => n2371, Z => 
                           n5264);
   U1506 : AO4 port map( A => n3072, B => n414, C => n371, D => n2370, Z => 
                           n5265);
   U1507 : AO4 port map( A => n3073, B => n415, C => n2448, D => n2369, Z => 
                           n5266);
   U1508 : AO4 port map( A => n3070, B => n416, C => n371, D => n2368, Z => 
                           n5267);
   U1509 : AO4 port map( A => n3071, B => n417, C => n371, D => n2367, Z => 
                           n5268);
   U1510 : AO4 port map( A => n3084, B => n418, C => n371, D => n2366, Z => 
                           n5269);
   U1511 : AO4 port map( A => n3085, B => n423, C => n371, D => n2365, Z => 
                           n5270);
   U1512 : AO4 port map( A => n3082, B => n424, C => n371, D => n2364, Z => 
                           n5271);
   U1513 : AO4 port map( A => n3083, B => n425, C => n371, D => n2363, Z => 
                           n5272);
   U1514 : AO4 port map( A => n3080, B => n426, C => n371, D => n2362, Z => 
                           n5273);
   U1515 : AO4 port map( A => n3081, B => n427, C => n371, D => n2361, Z => 
                           n5274);
   U1516 : AO4 port map( A => n3078, B => n428, C => n371, D => n2360, Z => 
                           n5275);
   U1517 : AO4 port map( A => n3079, B => n429, C => n371, D => n2359, Z => 
                           n5276);
   U1518 : AO4 port map( A => n3028, B => n751, C => n371, D => n2358, Z => 
                           n5277);
   U1519 : AO4 port map( A => n3029, B => n795, C => n371, D => n2357, Z => 
                           n5278);
   U1521 : AO4 port map( A => n3026, B => n839, C => n371, D => n2356, Z => 
                           n5279);
   U1522 : AO4 port map( A => n3027, B => n883, C => n371, D => n2355, Z => 
                           n5280);
   U1523 : AO4 port map( A => n3024, B => n430, C => n371, D => n2354, Z => 
                           n5281);
   U1524 : AO4 port map( A => n3025, B => n435, C => n371, D => n2353, Z => 
                           n5282);
   U1525 : AO4 port map( A => n3022, B => n436, C => n371, D => n2352, Z => 
                           n5283);
   U1526 : AO4 port map( A => n3023, B => n437, C => n371, D => n2351, Z => 
                           n5284);
   U1527 : AO4 port map( A => n3036, B => n927, C => n371, D => n2350, Z => 
                           n5285);
   U1528 : AO4 port map( A => n3037, B => n971, C => n371, D => n2349, Z => 
                           n5286);
   U1529 : AO4 port map( A => n3034, B => n1015, C => n371, D => n2348, Z => 
                           n5287);
   U1530 : AO4 port map( A => n3035, B => n1059, C => n371, D => n2347, Z => 
                           n5288);
   U1531 : AO4 port map( A => n3032, B => n438, C => n371, D => n2346, Z => 
                           n5289);
   U1532 : AO4 port map( A => n3033, B => n439, C => n371, D => n2345, Z => 
                           n5290);
   U1533 : AO4 port map( A => n3030, B => n440, C => n2448, D => n2344, Z => 
                           n5291);
   U1534 : AO4 port map( A => n3031, B => n441, C => n2448, D => n2343, Z => 
                           n5292);
   U1535 : AO4 port map( A => n3044, B => n1103, C => n2448, D => n2342, Z => 
                           n5293);
   U1536 : AO4 port map( A => n3045, B => n1147, C => n2448, D => n2341, Z => 
                           n5294);
   U1537 : AO4 port map( A => n3042, B => n1191, C => n2448, D => n2340, Z => 
                           n5295);
   U1538 : AO4 port map( A => n3043, B => n1235, C => n371, D => n2339, Z => 
                           n5296);
   U1539 : AO4 port map( A => n3040, B => n442, C => n2448, D => n2338, Z => 
                           n5297);
   U1540 : AO4 port map( A => n3041, B => n443, C => n2448, D => n2337, Z => 
                           n5298);
   U1541 : AO4 port map( A => n3038, B => n487, C => n371, D => n2336, Z => 
                           n5299);
   U1542 : AO4 port map( A => n3039, B => n531, C => n2448, D => n2335, Z => 
                           n5300);
   U1543 : AO4 port map( A => n3052, B => n1279, C => n2448, D => n2334, Z => 
                           n5301);
   U1544 : AO4 port map( A => n3053, B => n1323, C => n371, D => n2333, Z => 
                           n5302);
   U1545 : AO4 port map( A => n3050, B => n1367, C => n2448, D => n2332, Z => 
                           n5303);
   U1546 : AO4 port map( A => n3051, B => n1411, C => n2448, D => n2331, Z => 
                           n5304);
   U1547 : AO4 port map( A => n3048, B => n575, C => n371, D => n2330, Z => 
                           n5305);
   U1548 : AO4 port map( A => n3049, B => n619, C => n2448, D => n2329, Z => 
                           n5306);
   U1549 : AO4 port map( A => n3046, B => n663, C => n2448, D => n2328, Z => 
                           n5307);
   U1550 : AO4 port map( A => n3047, B => n707, C => n371, D => n2327, Z => 
                           n5308);
   U1551 : AO4 port map( A => n3132, B => n390, C => n349, D => n2382, Z => 
                           n5765);
   U1552 : AO4 port map( A => n3133, B => n399, C => n2456, D => n2381, Z => 
                           n5766);
   U1553 : AO4 port map( A => n3130, B => n400, C => n349, D => n2380, Z => 
                           n5767);
   U1554 : AO4 port map( A => n3131, B => n401, C => n2456, D => n2379, Z => 
                           n5768);
   U1555 : AO4 port map( A => n3128, B => n402, C => n349, D => n2378, Z => 
                           n5769);
   U1556 : AO4 port map( A => n3129, B => n403, C => n2456, D => n2377, Z => 
                           n5770);
   U1557 : AO4 port map( A => n3126, B => n404, C => n349, D => n2376, Z => 
                           n5771);
   U1558 : AO4 port map( A => n3127, B => n405, C => n2456, D => n2375, Z => 
                           n5772);
   U1559 : AO4 port map( A => n3140, B => n406, C => n349, D => n2374, Z => 
                           n5773);
   U1560 : AO4 port map( A => n3141, B => n411, C => n2456, D => n2373, Z => 
                           n5774);
   U1561 : AO4 port map( A => n3138, B => n412, C => n2456, D => n2372, Z => 
                           n5775);
   U1562 : AO4 port map( A => n3139, B => n413, C => n2456, D => n2371, Z => 
                           n5776);
   U1563 : AO4 port map( A => n3136, B => n414, C => n2456, D => n2370, Z => 
                           n5777);
   U1565 : AO4 port map( A => n3137, B => n415, C => n2456, D => n2369, Z => 
                           n5778);
   U1566 : AO4 port map( A => n3134, B => n416, C => n349, D => n2368, Z => 
                           n5779);
   U1567 : AO4 port map( A => n3135, B => n417, C => n2456, D => n2367, Z => 
                           n5780);
   U1568 : AO4 port map( A => n3148, B => n418, C => n2456, D => n2366, Z => 
                           n5781);
   U1569 : AO4 port map( A => n3149, B => n423, C => n349, D => n2365, Z => 
                           n5782);
   U1570 : AO4 port map( A => n3146, B => n424, C => n2456, D => n2364, Z => 
                           n5783);
   U1571 : AO4 port map( A => n3147, B => n425, C => n2456, D => n2363, Z => 
                           n5784);
   U1572 : AO4 port map( A => n3144, B => n426, C => n349, D => n2362, Z => 
                           n5785);
   U1573 : AO4 port map( A => n3145, B => n427, C => n2456, D => n2361, Z => 
                           n5786);
   U1574 : AO4 port map( A => n3142, B => n428, C => n2456, D => n2360, Z => 
                           n5787);
   U1575 : AO4 port map( A => n3143, B => n429, C => n349, D => n2359, Z => 
                           n5788);
   U1576 : AO4 port map( A => n3092, B => n751, C => n2456, D => n2358, Z => 
                           n5789);
   U1577 : AO4 port map( A => n3093, B => n795, C => n2456, D => n2357, Z => 
                           n5790);
   U1578 : AO4 port map( A => n3090, B => n839, C => n349, D => n2356, Z => 
                           n5791);
   U1579 : AO4 port map( A => n3091, B => n883, C => n2456, D => n2355, Z => 
                           n5792);
   U1580 : AO4 port map( A => n3088, B => n430, C => n349, D => n2354, Z => 
                           n5793);
   U1581 : AO4 port map( A => n3089, B => n435, C => n349, D => n2353, Z => 
                           n5794);
   U1582 : AO4 port map( A => n3086, B => n436, C => n349, D => n2352, Z => 
                           n5795);
   U1583 : AO4 port map( A => n3087, B => n437, C => n349, D => n2351, Z => 
                           n5796);
   U1584 : AO4 port map( A => n3100, B => n927, C => n349, D => n2350, Z => 
                           n5797);
   U1585 : AO4 port map( A => n3101, B => n971, C => n349, D => n2349, Z => 
                           n5798);
   U1586 : AO4 port map( A => n3098, B => n1015, C => n349, D => n2348, Z => 
                           n5799);
   U1587 : AO4 port map( A => n3099, B => n1059, C => n349, D => n2347, Z => 
                           n5800);
   U1588 : AO4 port map( A => n3096, B => n438, C => n349, D => n2346, Z => 
                           n5801);
   U1589 : AO4 port map( A => n3097, B => n439, C => n349, D => n2345, Z => 
                           n5802);
   U1590 : AO4 port map( A => n3094, B => n440, C => n349, D => n2344, Z => 
                           n5803);
   U1591 : AO4 port map( A => n3095, B => n441, C => n349, D => n2343, Z => 
                           n5804);
   U1592 : AO4 port map( A => n3108, B => n1103, C => n349, D => n2342, Z => 
                           n5805);
   U1593 : AO4 port map( A => n3109, B => n1147, C => n349, D => n2341, Z => 
                           n5806);
   U1594 : AO4 port map( A => n3106, B => n1191, C => n349, D => n2340, Z => 
                           n5807);
   U1595 : AO4 port map( A => n3107, B => n1235, C => n349, D => n2339, Z => 
                           n5808);
   U1596 : AO4 port map( A => n3104, B => n442, C => n349, D => n2338, Z => 
                           n5809);
   U1597 : AO4 port map( A => n3105, B => n443, C => n349, D => n2337, Z => 
                           n5810);
   U1598 : AO4 port map( A => n3102, B => n487, C => n349, D => n2336, Z => 
                           n5811);
   U1599 : AO4 port map( A => n3103, B => n531, C => n2456, D => n2335, Z => 
                           n5812);
   U1600 : AO4 port map( A => n3116, B => n1279, C => n2456, D => n2334, Z => 
                           n5813);
   U1601 : AO4 port map( A => n3117, B => n1323, C => n2456, D => n2333, Z => 
                           n5814);
   U1602 : AO4 port map( A => n3114, B => n1367, C => n2456, D => n2332, Z => 
                           n5815);
   U1603 : AO4 port map( A => n3115, B => n1411, C => n2456, D => n2331, Z => 
                           n5816);
   U1604 : AO4 port map( A => n3112, B => n575, C => n2456, D => n2330, Z => 
                           n5817);
   U1605 : AO4 port map( A => n3113, B => n619, C => n2456, D => n2329, Z => 
                           n5818);
   U1606 : AO4 port map( A => n3110, B => n663, C => n2456, D => n2328, Z => 
                           n5819);
   U1607 : AO4 port map( A => n3111, B => n707, C => n2456, D => n2327, Z => 
                           n5820);
   U1609 : AO4 port map( A => n3196, B => n390, C => n2464, D => n2382, Z => 
                           n6277);
   U1610 : AO4 port map( A => n3197, B => n399, C => n2464, D => n2381, Z => 
                           n6278);
   U1611 : AO4 port map( A => n3194, B => n400, C => n2464, D => n2380, Z => 
                           n6279);
   U1612 : AO4 port map( A => n3195, B => n401, C => n2464, D => n2379, Z => 
                           n6280);
   U1613 : AO4 port map( A => n3192, B => n402, C => n2464, D => n2378, Z => 
                           n6281);
   U1614 : AO4 port map( A => n3193, B => n403, C => n2464, D => n2377, Z => 
                           n6282);
   U1615 : AO4 port map( A => n3190, B => n404, C => n2464, D => n2376, Z => 
                           n6283);
   U1616 : AO4 port map( A => n3191, B => n405, C => n2464, D => n2375, Z => 
                           n6284);
   U1617 : AO4 port map( A => n3204, B => n406, C => n348, D => n2374, Z => 
                           n6285);
   U1618 : AO4 port map( A => n3205, B => n411, C => n2464, D => n2373, Z => 
                           n6286);
   U1619 : AO4 port map( A => n3202, B => n412, C => n2464, D => n2372, Z => 
                           n6287);
   U1620 : AO4 port map( A => n3203, B => n413, C => n2464, D => n2371, Z => 
                           n6288);
   U1621 : AO4 port map( A => n3200, B => n414, C => n348, D => n2370, Z => 
                           n6289);
   U1622 : AO4 port map( A => n3201, B => n415, C => n2464, D => n2369, Z => 
                           n6290);
   U1623 : AO4 port map( A => n3198, B => n416, C => n348, D => n2368, Z => 
                           n6291);
   U1624 : AO4 port map( A => n3199, B => n417, C => n348, D => n2367, Z => 
                           n6292);
   U1625 : AO4 port map( A => n3212, B => n418, C => n348, D => n2366, Z => 
                           n6293);
   U1626 : AO4 port map( A => n3213, B => n423, C => n348, D => n2365, Z => 
                           n6294);
   U1627 : AO4 port map( A => n3210, B => n424, C => n348, D => n2364, Z => 
                           n6295);
   U1628 : AO4 port map( A => n3211, B => n425, C => n348, D => n2363, Z => 
                           n6296);
   U1629 : AO4 port map( A => n3208, B => n426, C => n348, D => n2362, Z => 
                           n6297);
   U1630 : AO4 port map( A => n3209, B => n427, C => n348, D => n2361, Z => 
                           n6298);
   U1631 : AO4 port map( A => n3206, B => n428, C => n348, D => n2360, Z => 
                           n6299);
   U1632 : AO4 port map( A => n3207, B => n429, C => n348, D => n2359, Z => 
                           n6300);
   U1633 : AO4 port map( A => n3156, B => n751, C => n348, D => n2358, Z => 
                           n6301);
   U1634 : AO4 port map( A => n3157, B => n795, C => n348, D => n2357, Z => 
                           n6302);
   U1635 : AO4 port map( A => n3154, B => n839, C => n348, D => n2356, Z => 
                           n6303);
   U1636 : AO4 port map( A => n3155, B => n883, C => n348, D => n2355, Z => 
                           n6304);
   U1637 : AO4 port map( A => n3152, B => n430, C => n348, D => n2354, Z => 
                           n6305);
   U1638 : AO4 port map( A => n3153, B => n435, C => n348, D => n2353, Z => 
                           n6306);
   U1639 : AO4 port map( A => n3150, B => n436, C => n348, D => n2352, Z => 
                           n6307);
   U1640 : AO4 port map( A => n3151, B => n437, C => n348, D => n2351, Z => 
                           n6308);
   U1641 : AO4 port map( A => n3164, B => n927, C => n348, D => n2350, Z => 
                           n6309);
   U1642 : AO4 port map( A => n3165, B => n971, C => n348, D => n2349, Z => 
                           n6310);
   U1643 : AO4 port map( A => n3162, B => n1015, C => n348, D => n2348, Z => 
                           n6311);
   U1644 : AO4 port map( A => n3163, B => n1059, C => n348, D => n2347, Z => 
                           n6312);
   U1645 : AO4 port map( A => n3160, B => n438, C => n348, D => n2346, Z => 
                           n6313);
   U1646 : AO4 port map( A => n3161, B => n439, C => n348, D => n2345, Z => 
                           n6314);
   U1647 : AO4 port map( A => n3158, B => n440, C => n2464, D => n2344, Z => 
                           n6315);
   U1648 : AO4 port map( A => n3159, B => n441, C => n2464, D => n2343, Z => 
                           n6316);
   U1649 : AO4 port map( A => n3172, B => n1103, C => n2464, D => n2342, Z => 
                           n6317);
   U1650 : AO4 port map( A => n3173, B => n1147, C => n2464, D => n2341, Z => 
                           n6318);
   U1651 : AO4 port map( A => n3170, B => n1191, C => n2464, D => n2340, Z => 
                           n6319);
   U1653 : AO4 port map( A => n3171, B => n1235, C => n348, D => n2339, Z => 
                           n6320);
   U1654 : AO4 port map( A => n3168, B => n442, C => n2464, D => n2338, Z => 
                           n6321);
   U1655 : AO4 port map( A => n3169, B => n443, C => n2464, D => n2337, Z => 
                           n6322);
   U1656 : AO4 port map( A => n3166, B => n487, C => n348, D => n2336, Z => 
                           n6323);
   U1657 : AO4 port map( A => n3167, B => n531, C => n2464, D => n2335, Z => 
                           n6324);
   U1658 : AO4 port map( A => n3180, B => n1279, C => n2464, D => n2334, Z => 
                           n6325);
   U1659 : AO4 port map( A => n3181, B => n1323, C => n348, D => n2333, Z => 
                           n6326);
   U1660 : AO4 port map( A => n3178, B => n1367, C => n2464, D => n2332, Z => 
                           n6327);
   U1661 : AO4 port map( A => n3179, B => n1411, C => n2464, D => n2331, Z => 
                           n6328);
   U1662 : AO4 port map( A => n3176, B => n575, C => n348, D => n2330, Z => 
                           n6329);
   U1663 : AO4 port map( A => n3177, B => n619, C => n2464, D => n2329, Z => 
                           n6330);
   U1664 : AO4 port map( A => n3174, B => n663, C => n2464, D => n2328, Z => 
                           n6331);
   U1665 : AO4 port map( A => n3175, B => n707, C => n348, D => n2327, Z => 
                           n6332);
   U1666 : AO4 port map( A => n3252, B => n378, C => n352, D => n2390, Z => 
                           n4733);
   U1667 : AO4 port map( A => n3253, B => n383, C => n2440, D => n2389, Z => 
                           n4734);
   U1668 : AO4 port map( A => n3250, B => n384, C => n2440, D => n2388, Z => 
                           n4735);
   U1669 : AO4 port map( A => n3251, B => n385, C => n2440, D => n2387, Z => 
                           n4736);
   U1670 : AO4 port map( A => n3248, B => n386, C => n352, D => n2386, Z => 
                           n4737);
   U1671 : AO4 port map( A => n3249, B => n387, C => n2440, D => n2385, Z => 
                           n4738);
   U1672 : AO4 port map( A => n3246, B => n388, C => n2440, D => n2384, Z => 
                           n4739);
   U1673 : AO4 port map( A => n3247, B => n389, C => n2440, D => n2383, Z => 
                           n4740);
   U1674 : AO4 port map( A => n3260, B => n390, C => n352, D => n2382, Z => 
                           n4741);
   U1675 : AO4 port map( A => n3261, B => n399, C => n2440, D => n2381, Z => 
                           n4742);
   U1676 : AO4 port map( A => n3258, B => n400, C => n352, D => n2380, Z => 
                           n4743);
   U1677 : AO4 port map( A => n3259, B => n401, C => n2440, D => n2379, Z => 
                           n4744);
   U1678 : AO4 port map( A => n3256, B => n402, C => n352, D => n2378, Z => 
                           n4745);
   U1679 : AO4 port map( A => n3257, B => n403, C => n2440, D => n2377, Z => 
                           n4746);
   U1680 : AO4 port map( A => n3254, B => n404, C => n352, D => n2376, Z => 
                           n4747);
   U1681 : AO4 port map( A => n3255, B => n405, C => n2440, D => n2375, Z => 
                           n4748);
   U1682 : AO4 port map( A => n3268, B => n406, C => n352, D => n2374, Z => 
                           n4749);
   U1683 : AO4 port map( A => n3269, B => n411, C => n2440, D => n2373, Z => 
                           n4750);
   U1684 : AO4 port map( A => n3266, B => n412, C => n2440, D => n2372, Z => 
                           n4751);
   U1685 : AO4 port map( A => n3267, B => n413, C => n2440, D => n2371, Z => 
                           n4752);
   U1686 : AO4 port map( A => n3264, B => n414, C => n2440, D => n2370, Z => 
                           n4753);
   U1687 : AO4 port map( A => n3265, B => n415, C => n2440, D => n2369, Z => 
                           n4754);
   U1688 : AO4 port map( A => n3262, B => n416, C => n352, D => n2368, Z => 
                           n4755);
   U1689 : AO4 port map( A => n3263, B => n417, C => n2440, D => n2367, Z => 
                           n4756);
   U1690 : AO4 port map( A => n3276, B => n418, C => n2440, D => n2366, Z => 
                           n4757);
   U1691 : AO4 port map( A => n3277, B => n423, C => n352, D => n2365, Z => 
                           n4758);
   U1692 : AO4 port map( A => n3274, B => n424, C => n2440, D => n2364, Z => 
                           n4759);
   U1693 : AO4 port map( A => n3275, B => n425, C => n2440, D => n2363, Z => 
                           n4760);
   U1694 : AO4 port map( A => n3272, B => n426, C => n352, D => n2362, Z => 
                           n4761);
   U1695 : AO4 port map( A => n3273, B => n427, C => n2440, D => n2361, Z => 
                           n4762);
   U1697 : AO4 port map( A => n3270, B => n428, C => n2440, D => n2360, Z => 
                           n4763);
   U1698 : AO4 port map( A => n3271, B => n429, C => n352, D => n2359, Z => 
                           n4764);
   U1699 : AO4 port map( A => n3220, B => n751, C => n2440, D => n2358, Z => 
                           n4765);
   U1700 : AO4 port map( A => n3221, B => n795, C => n2440, D => n2357, Z => 
                           n4766);
   U1701 : AO4 port map( A => n3218, B => n839, C => n352, D => n2356, Z => 
                           n4767);
   U1702 : AO4 port map( A => n3219, B => n883, C => n2440, D => n2355, Z => 
                           n4768);
   U1703 : AO4 port map( A => n3216, B => n430, C => n352, D => n2354, Z => 
                           n4769);
   U1704 : AO4 port map( A => n3217, B => n435, C => n352, D => n2353, Z => 
                           n4770);
   U1705 : AO4 port map( A => n3214, B => n436, C => n352, D => n2352, Z => 
                           n4771);
   U1706 : AO4 port map( A => n3215, B => n437, C => n352, D => n2351, Z => 
                           n4772);
   U1707 : AO4 port map( A => n3228, B => n927, C => n352, D => n2350, Z => 
                           n4773);
   U1708 : AO4 port map( A => n3229, B => n971, C => n352, D => n2349, Z => 
                           n4774);
   U1709 : AO4 port map( A => n3226, B => n1015, C => n352, D => n2348, Z => 
                           n4775);
   U1710 : AO4 port map( A => n3227, B => n1059, C => n352, D => n2347, Z => 
                           n4776);
   U1711 : AO4 port map( A => n3224, B => n438, C => n352, D => n2346, Z => 
                           n4777);
   U1712 : AO4 port map( A => n3225, B => n439, C => n352, D => n2345, Z => 
                           n4778);
   U1713 : AO4 port map( A => n3222, B => n440, C => n352, D => n2344, Z => 
                           n4779);
   U1714 : AO4 port map( A => n3223, B => n441, C => n352, D => n2343, Z => 
                           n4780);
   U1715 : AO4 port map( A => n3236, B => n1103, C => n352, D => n2342, Z => 
                           n4781);
   U1716 : AO4 port map( A => n3237, B => n1147, C => n352, D => n2341, Z => 
                           n4782);
   U1717 : AO4 port map( A => n3234, B => n1191, C => n352, D => n2340, Z => 
                           n4783);
   U1718 : AO4 port map( A => n3235, B => n1235, C => n352, D => n2339, Z => 
                           n4784);
   U1719 : AO4 port map( A => n3232, B => n442, C => n352, D => n2338, Z => 
                           n4785);
   U1720 : AO4 port map( A => n3233, B => n443, C => n352, D => n2337, Z => 
                           n4786);
   U1721 : AO4 port map( A => n3230, B => n487, C => n352, D => n2336, Z => 
                           n4787);
   U1722 : AO4 port map( A => n3231, B => n531, C => n2440, D => n2335, Z => 
                           n4788);
   U1723 : AO4 port map( A => n3244, B => n1279, C => n2440, D => n2334, Z => 
                           n4789);
   U1724 : AO4 port map( A => n3245, B => n1323, C => n2440, D => n2333, Z => 
                           n4790);
   U1725 : AO4 port map( A => n3242, B => n1367, C => n2440, D => n2332, Z => 
                           n4791);
   U1726 : AO4 port map( A => n3243, B => n1411, C => n2440, D => n2331, Z => 
                           n4792);
   U1727 : AO4 port map( A => n3240, B => n575, C => n2440, D => n2330, Z => 
                           n4793);
   U1728 : AO4 port map( A => n3241, B => n619, C => n2440, D => n2329, Z => 
                           n4794);
   U1729 : AO4 port map( A => n3238, B => n663, C => n2440, D => n2328, Z => 
                           n4795);
   U1730 : AO4 port map( A => n3239, B => n707, C => n2440, D => n2327, Z => 
                           n4796);
   U1731 : AO4 port map( A => n3324, B => n390, C => n366, D => n2382, Z => 
                           n5317);
   U1732 : AO4 port map( A => n3325, B => n399, C => n2449, D => n2381, Z => 
                           n5318);
   U1733 : AO4 port map( A => n3322, B => n400, C => n366, D => n2380, Z => 
                           n5319);
   U1734 : AO4 port map( A => n3323, B => n401, C => n2449, D => n2379, Z => 
                           n5320);
   U1735 : AO4 port map( A => n3320, B => n402, C => n366, D => n2378, Z => 
                           n5321);
   U1736 : AO4 port map( A => n3321, B => n403, C => n2449, D => n2377, Z => 
                           n5322);
   U1737 : AO4 port map( A => n3318, B => n404, C => n366, D => n2376, Z => 
                           n5323);
   U1738 : AO4 port map( A => n3319, B => n405, C => n2449, D => n2375, Z => 
                           n5324);
   U1739 : AO4 port map( A => n3332, B => n406, C => n366, D => n2374, Z => 
                           n5325);
   U1741 : AO4 port map( A => n3333, B => n411, C => n2449, D => n2373, Z => 
                           n5326);
   U1742 : AO4 port map( A => n3330, B => n412, C => n2449, D => n2372, Z => 
                           n5327);
   U1743 : AO4 port map( A => n3331, B => n413, C => n2449, D => n2371, Z => 
                           n5328);
   U1744 : AO4 port map( A => n3328, B => n414, C => n2449, D => n2370, Z => 
                           n5329);
   U1745 : AO4 port map( A => n3329, B => n415, C => n2449, D => n2369, Z => 
                           n5330);
   U1746 : AO4 port map( A => n3326, B => n416, C => n366, D => n2368, Z => 
                           n5331);
   U1747 : AO4 port map( A => n3327, B => n417, C => n2449, D => n2367, Z => 
                           n5332);
   U1748 : AO4 port map( A => n3340, B => n418, C => n2449, D => n2366, Z => 
                           n5333);
   U1750 : AO4 port map( A => n3341, B => n423, C => n366, D => n2365, Z => 
                           n5334);
   U1751 : AO4 port map( A => n3338, B => n424, C => n2449, D => n2364, Z => 
                           n5335);
   U1752 : AO4 port map( A => n3339, B => n425, C => n2449, D => n2363, Z => 
                           n5336);
   U1753 : AO4 port map( A => n3336, B => n426, C => n366, D => n2362, Z => 
                           n5337);
   U1754 : AO4 port map( A => n3337, B => n427, C => n2449, D => n2361, Z => 
                           n5338);
   U1755 : AO4 port map( A => n3334, B => n428, C => n2449, D => n2360, Z => 
                           n5339);
   U1757 : AO4 port map( A => n3335, B => n429, C => n366, D => n2359, Z => 
                           n5340);
   U1758 : AO4 port map( A => n3284, B => n751, C => n2449, D => n2358, Z => 
                           n5341);
   U1759 : AO4 port map( A => n3285, B => n795, C => n2449, D => n2357, Z => 
                           n5342);
   U1760 : AO4 port map( A => n3282, B => n839, C => n366, D => n2356, Z => 
                           n5343);
   U1761 : AO4 port map( A => n3283, B => n883, C => n2449, D => n2355, Z => 
                           n5344);
   U1762 : AO4 port map( A => n3280, B => n430, C => n366, D => n2354, Z => 
                           n5345);
   U1763 : AO4 port map( A => n3281, B => n435, C => n366, D => n2353, Z => 
                           n5346);
   U1765 : AO4 port map( A => n3278, B => n436, C => n366, D => n2352, Z => 
                           n5347);
   U1766 : AO4 port map( A => n3279, B => n437, C => n366, D => n2351, Z => 
                           n5348);
   U1767 : AO4 port map( A => n3292, B => n927, C => n366, D => n2350, Z => 
                           n5349);
   U1768 : AO4 port map( A => n3293, B => n971, C => n366, D => n2349, Z => 
                           n5350);
   U1769 : AO4 port map( A => n3290, B => n1015, C => n366, D => n2348, Z => 
                           n5351);
   U1770 : AO4 port map( A => n3291, B => n1059, C => n366, D => n2347, Z => 
                           n5352);
   U1773 : AO4 port map( A => n3288, B => n438, C => n366, D => n2346, Z => 
                           n5353);
   U1774 : AO4 port map( A => n3289, B => n439, C => n366, D => n2345, Z => 
                           n5354);
   U1775 : AO4 port map( A => n3286, B => n440, C => n366, D => n2344, Z => 
                           n5355);
   U1776 : AO4 port map( A => n3287, B => n441, C => n366, D => n2343, Z => 
                           n5356);
   U1777 : AO4 port map( A => n3300, B => n1103, C => n366, D => n2342, Z => 
                           n5357);
   U1778 : AO4 port map( A => n3301, B => n1147, C => n366, D => n2341, Z => 
                           n5358);
   U1779 : AO4 port map( A => n3298, B => n1191, C => n366, D => n2340, Z => 
                           n5359);
   U1781 : AO4 port map( A => n3299, B => n1235, C => n366, D => n2339, Z => 
                           n5360);
   U1782 : AO4 port map( A => n3296, B => n442, C => n366, D => n2338, Z => 
                           n5361);
   U1783 : AO4 port map( A => n3297, B => n443, C => n366, D => n2337, Z => 
                           n5362);
   U1784 : AO4 port map( A => n3294, B => n487, C => n366, D => n2336, Z => 
                           n5363);
   U1785 : AO4 port map( A => n3295, B => n531, C => n2449, D => n2335, Z => 
                           n5364);
   U1786 : AO4 port map( A => n3308, B => n1279, C => n2449, D => n2334, Z => 
                           n5365);
   U1788 : AO4 port map( A => n3309, B => n1323, C => n2449, D => n2333, Z => 
                           n5366);
   U1789 : AO4 port map( A => n3306, B => n1367, C => n2449, D => n2332, Z => 
                           n5367);
   U1790 : AO4 port map( A => n3307, B => n1411, C => n2449, D => n2331, Z => 
                           n5368);
   U1791 : AO4 port map( A => n3304, B => n575, C => n2449, D => n2330, Z => 
                           n5369);
   U1792 : AO4 port map( A => n3305, B => n619, C => n2449, D => n2329, Z => 
                           n5370);
   U1793 : AO4 port map( A => n3302, B => n663, C => n2449, D => n2328, Z => 
                           n5371);
   U1794 : AO4 port map( A => n3303, B => n707, C => n2449, D => n2327, Z => 
                           n5372);
   U1796 : AO4 port map( A => n3388, B => n390, C => n347, D => n2382, Z => 
                           n5829);
   U1797 : AO4 port map( A => n3389, B => n399, C => n2457, D => n2381, Z => 
                           n5830);
   U1798 : AO4 port map( A => n3386, B => n400, C => n347, D => n2380, Z => 
                           n5831);
   U1799 : AO4 port map( A => n3387, B => n401, C => n2457, D => n2379, Z => 
                           n5832);
   U1800 : AO4 port map( A => n3384, B => n402, C => n347, D => n2378, Z => 
                           n5833);
   U1801 : AO4 port map( A => n3385, B => n403, C => n2457, D => n2377, Z => 
                           n5834);
   U1804 : AO4 port map( A => n3382, B => n404, C => n347, D => n2376, Z => 
                           n5835);
   U1805 : AO4 port map( A => n3383, B => n405, C => n2457, D => n2375, Z => 
                           n5836);
   U1806 : AO4 port map( A => n3396, B => n406, C => n347, D => n2374, Z => 
                           n5837);
   U1807 : AO4 port map( A => n3397, B => n411, C => n2457, D => n2373, Z => 
                           n5838);
   U1808 : AO4 port map( A => n3394, B => n412, C => n2457, D => n2372, Z => 
                           n5839);
   U1809 : AO4 port map( A => n3395, B => n413, C => n2457, D => n2371, Z => 
                           n5840);
   U1810 : AO4 port map( A => n3392, B => n414, C => n2457, D => n2370, Z => 
                           n5841);
   U1811 : AO4 port map( A => n3393, B => n415, C => n2457, D => n2369, Z => 
                           n5842);
   U1812 : AO4 port map( A => n3390, B => n416, C => n347, D => n2368, Z => 
                           n5843);
   U1814 : AO4 port map( A => n3391, B => n417, C => n2457, D => n2367, Z => 
                           n5844);
   U1815 : AO4 port map( A => n3404, B => n418, C => n2457, D => n2366, Z => 
                           n5845);
   U1816 : AO4 port map( A => n3405, B => n423, C => n347, D => n2365, Z => 
                           n5846);
   U1817 : AO4 port map( A => n3402, B => n424, C => n2457, D => n2364, Z => 
                           n5847);
   U1818 : AO4 port map( A => n3403, B => n425, C => n2457, D => n2363, Z => 
                           n5848);
   U1819 : AO4 port map( A => n3400, B => n426, C => n347, D => n2362, Z => 
                           n5849);
   U1821 : AO4 port map( A => n3401, B => n427, C => n2457, D => n2361, Z => 
                           n5850);
   U1822 : AO4 port map( A => n3398, B => n428, C => n2457, D => n2360, Z => 
                           n5851);
   U1823 : AO4 port map( A => n3399, B => n429, C => n347, D => n2359, Z => 
                           n5852);
   U1824 : AO4 port map( A => n3348, B => n751, C => n2457, D => n2358, Z => 
                           n5853);
   U1825 : AO4 port map( A => n3349, B => n795, C => n2457, D => n2357, Z => 
                           n5854);
   U1826 : AO4 port map( A => n3346, B => n839, C => n347, D => n2356, Z => 
                           n5855);
   U1827 : AO4 port map( A => n3347, B => n883, C => n2457, D => n2355, Z => 
                           n5856);
   U1829 : AO4 port map( A => n3344, B => n430, C => n347, D => n2354, Z => 
                           n5857);
   U1830 : AO4 port map( A => n3345, B => n435, C => n347, D => n2353, Z => 
                           n5858);
   U1831 : AO4 port map( A => n3342, B => n436, C => n347, D => n2352, Z => 
                           n5859);
   U1832 : AO4 port map( A => n3343, B => n437, C => n347, D => n2351, Z => 
                           n5860);
   U1833 : AO4 port map( A => n3356, B => n927, C => n347, D => n2350, Z => 
                           n5861);
   U1834 : AO4 port map( A => n3357, B => n971, C => n347, D => n2349, Z => 
                           n5862);
   U1837 : AO4 port map( A => n3354, B => n1015, C => n347, D => n2348, Z => 
                           n5863);
   U1838 : AO4 port map( A => n3355, B => n1059, C => n347, D => n2347, Z => 
                           n5864);
   U1839 : AO4 port map( A => n3352, B => n438, C => n347, D => n2346, Z => 
                           n5865);
   U1840 : AO4 port map( A => n3353, B => n439, C => n347, D => n2345, Z => 
                           n5866);
   U1841 : AO4 port map( A => n3350, B => n440, C => n347, D => n2344, Z => 
                           n5867);
   U1842 : AO4 port map( A => n3351, B => n441, C => n347, D => n2343, Z => 
                           n5868);
   U1843 : AO4 port map( A => n3364, B => n1103, C => n347, D => n2342, Z => 
                           n5869);
   U1844 : AO4 port map( A => n3365, B => n1147, C => n347, D => n2341, Z => 
                           n5870);
   U1847 : AO4 port map( A => n3362, B => n1191, C => n347, D => n2340, Z => 
                           n5871);
   U1848 : AO4 port map( A => n3363, B => n1235, C => n347, D => n2339, Z => 
                           n5872);
   U1849 : AO4 port map( A => n3360, B => n442, C => n347, D => n2338, Z => 
                           n5873);
   U1850 : AO4 port map( A => n3361, B => n443, C => n347, D => n2337, Z => 
                           n5874);
   U1851 : AO4 port map( A => n3358, B => n487, C => n347, D => n2336, Z => 
                           n5875);
   U1852 : AO4 port map( A => n3359, B => n531, C => n2457, D => n2335, Z => 
                           n5876);
   U1855 : AO4 port map( A => n3372, B => n1279, C => n2457, D => n2334, Z => 
                           n5877);
   U1856 : AO4 port map( A => n3373, B => n1323, C => n2457, D => n2333, Z => 
                           n5878);
   U1857 : AO4 port map( A => n3370, B => n1367, C => n2457, D => n2332, Z => 
                           n5879);
   U1858 : AO4 port map( A => n3371, B => n1411, C => n2457, D => n2331, Z => 
                           n5880);
   U1859 : AO4 port map( A => n3368, B => n575, C => n2457, D => n2330, Z => 
                           n5881);
   U1860 : AO4 port map( A => n3369, B => n619, C => n2457, D => n2329, Z => 
                           n5882);
   U1861 : AO4 port map( A => n3366, B => n663, C => n2457, D => n2328, Z => 
                           n5883);
   U1862 : AO4 port map( A => n3367, B => n707, C => n2457, D => n2327, Z => 
                           n5884);
   U1865 : AO4 port map( A => n3452, B => n390, C => n335, D => n2382, Z => 
                           n6341);
   U1866 : AO4 port map( A => n3453, B => n399, C => n335, D => n2381, Z => 
                           n6342);
   U1867 : AO4 port map( A => n3450, B => n400, C => n335, D => n2380, Z => 
                           n6343);
   U1869 : AO4 port map( A => n3451, B => n401, C => n2465, D => n2379, Z => 
                           n6344);
   U1871 : AO4 port map( A => n3448, B => n402, C => n2465, D => n2378, Z => 
                           n6345);
   U1872 : AO4 port map( A => n3449, B => n403, C => n2465, D => n2377, Z => 
                           n6346);
   U1873 : AO4 port map( A => n3446, B => n404, C => n2465, D => n2376, Z => 
                           n6347);
   U1875 : AO4 port map( A => n3447, B => n405, C => n2465, D => n2375, Z => 
                           n6348);
   U1876 : AO4 port map( A => n3460, B => n406, C => n2465, D => n2374, Z => 
                           n6349);
   U1878 : AO4 port map( A => n3461, B => n411, C => n2465, D => n2373, Z => 
                           n6350);
   U1879 : AO4 port map( A => n3458, B => n412, C => n2465, D => n2372, Z => 
                           n6351);
   U1882 : AO4 port map( A => n3459, B => n413, C => n2465, D => n2371, Z => 
                           n6352);
   U1883 : AO4 port map( A => n3456, B => n414, C => n2465, D => n2370, Z => 
                           n6353);
   U1885 : AO4 port map( A => n3457, B => n415, C => n2465, D => n2369, Z => 
                           n6354);
   U1886 : AO4 port map( A => n3454, B => n416, C => n335, D => n2368, Z => 
                           n6355);
   U1887 : AO4 port map( A => n3455, B => n417, C => n2465, D => n2367, Z => 
                           n6356);
   U1888 : AO4 port map( A => n3468, B => n418, C => n335, D => n2366, Z => 
                           n6357);
   U1890 : AO4 port map( A => n3469, B => n423, C => n2465, D => n2365, Z => 
                           n6358);
   U1891 : AO4 port map( A => n3466, B => n424, C => n335, D => n2364, Z => 
                           n6359);
   U1894 : AO4 port map( A => n3467, B => n425, C => n2465, D => n2363, Z => 
                           n6360);
   U1895 : AO4 port map( A => n3464, B => n426, C => n335, D => n2362, Z => 
                           n6361);
   U1898 : AO4 port map( A => n3465, B => n427, C => n2465, D => n2361, Z => 
                           n6362);
   U1899 : AO4 port map( A => n3462, B => n428, C => n2465, D => n2360, Z => 
                           n6363);
   U1900 : AO4 port map( A => n3463, B => n429, C => n2465, D => n2359, Z => 
                           n6364);
   U1901 : AO4 port map( A => n3412, B => n751, C => n2465, D => n2358, Z => 
                           n6365);
   U1902 : AO4 port map( A => n3413, B => n795, C => n2465, D => n2357, Z => 
                           n6366);
   U1903 : AO4 port map( A => n3410, B => n839, C => n2465, D => n2356, Z => 
                           n6367);
   U1904 : AO4 port map( A => n3411, B => n883, C => n2465, D => n2355, Z => 
                           n6368);
   U1905 : AO4 port map( A => n3408, B => n430, C => n335, D => n2354, Z => 
                           n6369);
   U1908 : AO4 port map( A => n3409, B => n435, C => n2465, D => n2353, Z => 
                           n6370);
   U1909 : AO4 port map( A => n3406, B => n436, C => n2465, D => n2352, Z => 
                           n6371);
   U1910 : AO4 port map( A => n3407, B => n437, C => n335, D => n2351, Z => 
                           n6372);
   U1912 : AO4 port map( A => n3420, B => n927, C => n2465, D => n2350, Z => 
                           n6373);
   U1913 : AO4 port map( A => n3421, B => n971, C => n2465, D => n2349, Z => 
                           n6374);
   U1916 : AO4 port map( A => n3418, B => n1015, C => n335, D => n2348, Z => 
                           n6375);
   U1918 : AO4 port map( A => n3419, B => n1059, C => n335, D => n2347, Z => 
                           n6376);
   U1919 : AO4 port map( A => n3416, B => n438, C => n335, D => n2346, Z => 
                           n6377);
   U1920 : AO4 port map( A => n3417, B => n439, C => n335, D => n2345, Z => 
                           n6378);
   U1921 : AO4 port map( A => n3414, B => n440, C => n335, D => n2344, Z => 
                           n6379);
   U1922 : AO4 port map( A => n3415, B => n441, C => n335, D => n2343, Z => 
                           n6380);
   U1923 : AO4 port map( A => n3428, B => n1103, C => n2465, D => n2342, Z => 
                           n6381);
   U1924 : AO4 port map( A => n3429, B => n1147, C => n2465, D => n2341, Z => 
                           n6382);
   U1925 : AO4 port map( A => n3426, B => n1191, C => n335, D => n2340, Z => 
                           n6383);
   U1926 : AO4 port map( A => n3427, B => n1235, C => n335, D => n2339, Z => 
                           n6384);
   U1927 : AO4 port map( A => n3424, B => n442, C => n335, D => n2338, Z => 
                           n6385);
   U1929 : AO4 port map( A => n3425, B => n443, C => n335, D => n2337, Z => 
                           n6386);
   U1930 : AO4 port map( A => n3422, B => n487, C => n335, D => n2336, Z => 
                           n6387);
   U1932 : AO4 port map( A => n3423, B => n531, C => n335, D => n2335, Z => 
                           n6388);
   U1933 : AO4 port map( A => n3436, B => n1279, C => n335, D => n2334, Z => 
                           n6389);
   U1934 : AO4 port map( A => n3437, B => n1323, C => n335, D => n2333, Z => 
                           n6390);
   U1935 : AO4 port map( A => n3434, B => n1367, C => n335, D => n2332, Z => 
                           n6391);
   U1936 : AO4 port map( A => n3435, B => n1411, C => n335, D => n2331, Z => 
                           n6392);
   U1937 : AO4 port map( A => n3432, B => n575, C => n335, D => n2330, Z => 
                           n6393);
   U1938 : AO4 port map( A => n3433, B => n619, C => n335, D => n2329, Z => 
                           n6394);
   U1939 : AO4 port map( A => n3430, B => n663, C => n335, D => n2328, Z => 
                           n6395);
   U1942 : AO4 port map( A => n3431, B => n707, C => n335, D => n2327, Z => 
                           n6396);
   U1944 : AO4 port map( A => n3508, B => n378, C => n2441, D => n2390, Z => 
                           n4797);
   U1945 : AO4 port map( A => n3509, B => n383, C => n2441, D => n2389, Z => 
                           n4798);
   U1949 : AO4 port map( A => n3506, B => n384, C => n2441, D => n2388, Z => 
                           n4799);
   U1950 : AO4 port map( A => n3507, B => n385, C => n2441, D => n2387, Z => 
                           n4800);
   U1951 : AO4 port map( A => n3504, B => n386, C => n2441, D => n2386, Z => 
                           n4801);
   U1953 : AO4 port map( A => n3505, B => n387, C => n2441, D => n2385, Z => 
                           n4802);
   U1954 : AO4 port map( A => n3502, B => n388, C => n2441, D => n2384, Z => 
                           n4803);
   U1955 : AO4 port map( A => n3503, B => n389, C => n2441, D => n2383, Z => 
                           n4804);
   U1957 : AO4 port map( A => n3516, B => n390, C => n2441, D => n2382, Z => 
                           n4805);
   U1959 : AO4 port map( A => n3517, B => n399, C => n2441, D => n2381, Z => 
                           n4806);
   U1960 : AO4 port map( A => n3514, B => n400, C => n2441, D => n2380, Z => 
                           n4807);
   U1962 : AO4 port map( A => n3515, B => n401, C => n2441, D => n2379, Z => 
                           n4808);
   U1963 : AO4 port map( A => n3512, B => n402, C => n2441, D => n2378, Z => 
                           n4809);
   U1964 : AO4 port map( A => n3513, B => n403, C => n2441, D => n2377, Z => 
                           n4810);
   U1965 : AO4 port map( A => n3510, B => n404, C => n2441, D => n2376, Z => 
                           n4811);
   U1966 : AO4 port map( A => n3511, B => n405, C => n2441, D => n2375, Z => 
                           n4812);
   U1967 : AO4 port map( A => n3524, B => n406, C => n376, D => n2374, Z => 
                           n4813);
   U1968 : AO4 port map( A => n3525, B => n411, C => n2441, D => n2373, Z => 
                           n4814);
   U1969 : AO4 port map( A => n3522, B => n412, C => n2441, D => n2372, Z => 
                           n4815);
   U1970 : AO4 port map( A => n3523, B => n413, C => n2441, D => n2371, Z => 
                           n4816);
   U1971 : AO4 port map( A => n3520, B => n414, C => n376, D => n2370, Z => 
                           n4817);
   U1972 : AO4 port map( A => n3521, B => n415, C => n2441, D => n2369, Z => 
                           n4818);
   U1973 : AO4 port map( A => n3518, B => n416, C => n376, D => n2368, Z => 
                           n4819);
   U1974 : AO4 port map( A => n3519, B => n417, C => n376, D => n2367, Z => 
                           n4820);
   U1976 : AO4 port map( A => n3532, B => n418, C => n376, D => n2366, Z => 
                           n4821);
   U1977 : AO4 port map( A => n3533, B => n423, C => n376, D => n2365, Z => 
                           n4822);
   U1978 : AO4 port map( A => n3530, B => n424, C => n376, D => n2364, Z => 
                           n4823);
   U1979 : AO4 port map( A => n3531, B => n425, C => n376, D => n2363, Z => 
                           n4824);
   U1980 : AO4 port map( A => n3528, B => n426, C => n376, D => n2362, Z => 
                           n4825);
   U1981 : AO4 port map( A => n3529, B => n427, C => n376, D => n2361, Z => 
                           n4826);
   U1985 : AO4 port map( A => n3526, B => n428, C => n376, D => n2360, Z => 
                           n4827);
   U1986 : AO4 port map( A => n3527, B => n429, C => n376, D => n2359, Z => 
                           n4828);
   U1987 : AO4 port map( A => n3476, B => n751, C => n376, D => n2358, Z => 
                           n4829);
   U1988 : AO4 port map( A => n3477, B => n795, C => n376, D => n2357, Z => 
                           n4830);
   U1990 : AO4 port map( A => n3474, B => n839, C => n376, D => n2356, Z => 
                           n4831);
   U1991 : AO4 port map( A => n3475, B => n883, C => n376, D => n2355, Z => 
                           n4832);
   U1993 : AO4 port map( A => n3472, B => n430, C => n376, D => n2354, Z => 
                           n4833);
   U1996 : AO4 port map( A => n3473, B => n435, C => n376, D => n2353, Z => 
                           n4834);
   U1997 : AO4 port map( A => n3470, B => n436, C => n376, D => n2352, Z => 
                           n4835);
   U1998 : AO4 port map( A => n3471, B => n437, C => n376, D => n2351, Z => 
                           n4836);
   U1999 : AO4 port map( A => n3484, B => n927, C => n376, D => n2350, Z => 
                           n4837);
   U2000 : AO4 port map( A => n3485, B => n971, C => n376, D => n2349, Z => 
                           n4838);
   U2001 : AO4 port map( A => n3482, B => n1015, C => n376, D => n2348, Z => 
                           n4839);
   U2002 : AO4 port map( A => n3483, B => n1059, C => n376, D => n2347, Z => 
                           n4840);
   U2003 : AO4 port map( A => n3480, B => n438, C => n376, D => n2346, Z => 
                           n4841);
   U2006 : AO4 port map( A => n3481, B => n439, C => n376, D => n2345, Z => 
                           n4842);
   U2007 : AO4 port map( A => n3478, B => n440, C => n2441, D => n2344, Z => 
                           n4843);
   U2008 : AO4 port map( A => n3479, B => n441, C => n2441, D => n2343, Z => 
                           n4844);
   U2009 : AO4 port map( A => n3492, B => n1103, C => n2441, D => n2342, Z => 
                           n4845);
   U2010 : AO4 port map( A => n3493, B => n1147, C => n2441, D => n2341, Z => 
                           n4846);
   U2012 : AO4 port map( A => n3490, B => n1191, C => n2441, D => n2340, Z => 
                           n4847);
   U2014 : AO4 port map( A => n3491, B => n1235, C => n376, D => n2339, Z => 
                           n4848);
   U2015 : AO4 port map( A => n3488, B => n442, C => n2441, D => n2338, Z => 
                           n4849);
   U2016 : AO4 port map( A => n3489, B => n443, C => n2441, D => n2337, Z => 
                           n4850);
   U2017 : AO4 port map( A => n3486, B => n487, C => n376, D => n2336, Z => 
                           n4851);
   U2018 : AO4 port map( A => n3487, B => n531, C => n2441, D => n2335, Z => 
                           n4852);
   U2020 : AO4 port map( A => n3500, B => n1279, C => n2441, D => n2334, Z => 
                           n4853);
   U2021 : AO4 port map( A => n3501, B => n1323, C => n376, D => n2333, Z => 
                           n4854);
   U2022 : AO4 port map( A => n3498, B => n1367, C => n2441, D => n2332, Z => 
                           n4855);
   U2023 : AO4 port map( A => n3499, B => n1411, C => n2441, D => n2331, Z => 
                           n4856);
   U2024 : AO4 port map( A => n3496, B => n575, C => n376, D => n2330, Z => 
                           n4857);
   U2025 : AO4 port map( A => n3497, B => n619, C => n2441, D => n2329, Z => 
                           n4858);
   U2027 : AO4 port map( A => n3494, B => n663, C => n2441, D => n2328, Z => 
                           n4859);
   U2029 : AO4 port map( A => n3495, B => n707, C => n376, D => n2327, Z => 
                           n4860);
   U2030 : AO4 port map( A => n3580, B => n390, C => n365, D => n2382, Z => 
                           n5381);
   U2031 : AO4 port map( A => n3581, B => n399, C => n365, D => n2381, Z => 
                           n5382);
   U2032 : AO4 port map( A => n3578, B => n400, C => n365, D => n2380, Z => 
                           n5383);
   U2034 : AO4 port map( A => n3579, B => n401, C => n2450, D => n2379, Z => 
                           n5384);
   U2036 : AO4 port map( A => n3576, B => n402, C => n2450, D => n2378, Z => 
                           n5385);
   U2038 : AO4 port map( A => n3577, B => n403, C => n2450, D => n2377, Z => 
                           n5386);
   U2039 : AO4 port map( A => n3574, B => n404, C => n2450, D => n2376, Z => 
                           n5387);
   U2040 : AO4 port map( A => n3575, B => n405, C => n2450, D => n2375, Z => 
                           n5388);
   U2041 : AO4 port map( A => n3588, B => n406, C => n2450, D => n2374, Z => 
                           n5389);
   U2042 : AO4 port map( A => n3589, B => n411, C => n2450, D => n2373, Z => 
                           n5390);
   U2044 : AO4 port map( A => n3586, B => n412, C => n2450, D => n2372, Z => 
                           n5391);
   U2045 : AO4 port map( A => n3587, B => n413, C => n2450, D => n2371, Z => 
                           n5392);
   U2046 : AO4 port map( A => n3584, B => n414, C => n2450, D => n2370, Z => 
                           n5393);
   U2047 : AO4 port map( A => n3585, B => n415, C => n2450, D => n2369, Z => 
                           n5394);
   U2049 : AO4 port map( A => n3582, B => n416, C => n365, D => n2368, Z => 
                           n5395);
   U2050 : AO4 port map( A => n3583, B => n417, C => n2450, D => n2367, Z => 
                           n5396);
   U2052 : AO4 port map( A => n3596, B => n418, C => n365, D => n2366, Z => 
                           n5397);
   U2053 : AO4 port map( A => n3597, B => n423, C => n2450, D => n2365, Z => 
                           n5398);
   U2054 : AO4 port map( A => n3594, B => n424, C => n365, D => n2364, Z => 
                           n5399);
   U2055 : AO4 port map( A => n3595, B => n425, C => n2450, D => n2363, Z => 
                           n5400);
   U2056 : AO4 port map( A => n3592, B => n426, C => n365, D => n2362, Z => 
                           n5401);
   U2057 : AO4 port map( A => n3593, B => n427, C => n2450, D => n2361, Z => 
                           n5402);
   U2058 : AO4 port map( A => n3590, B => n428, C => n2450, D => n2360, Z => 
                           n5403);
   U2059 : AO4 port map( A => n3591, B => n429, C => n2450, D => n2359, Z => 
                           n5404);
   U2060 : AO4 port map( A => n3540, B => n751, C => n2450, D => n2358, Z => 
                           n5405);
   U2061 : AO4 port map( A => n3541, B => n795, C => n2450, D => n2357, Z => 
                           n5406);
   U2062 : AO4 port map( A => n3538, B => n839, C => n2450, D => n2356, Z => 
                           n5407);
   U2063 : AO4 port map( A => n3539, B => n883, C => n2450, D => n2355, Z => 
                           n5408);
   U2064 : AO4 port map( A => n3536, B => n430, C => n365, D => n2354, Z => 
                           n5409);
   U2066 : AO4 port map( A => n3537, B => n435, C => n2450, D => n2353, Z => 
                           n5410);
   U2067 : AO4 port map( A => n3534, B => n436, C => n2450, D => n2352, Z => 
                           n5411);
   U2068 : AO4 port map( A => n3535, B => n437, C => n365, D => n2351, Z => 
                           n5412);
   U2069 : AO4 port map( A => n3548, B => n927, C => n2450, D => n2350, Z => 
                           n5413);
   U2070 : AO4 port map( A => n3549, B => n971, C => n2450, D => n2349, Z => 
                           n5414);
   U2071 : AO4 port map( A => n3546, B => n1015, C => n365, D => n2348, Z => 
                           n5415);
   U2073 : AO4 port map( A => n3547, B => n1059, C => n365, D => n2347, Z => 
                           n5416);
   U2078 : AO4 port map( A => n3544, B => n438, C => n365, D => n2346, Z => 
                           n5417);
   U2079 : AO4 port map( A => n3545, B => n439, C => n365, D => n2345, Z => 
                           n5418);
   U2080 : AO4 port map( A => n3542, B => n440, C => n365, D => n2344, Z => 
                           n5419);
   U2082 : AO4 port map( A => n3543, B => n441, C => n365, D => n2343, Z => 
                           n5420);
   U2083 : AO4 port map( A => n3556, B => n1103, C => n2450, D => n2342, Z => 
                           n5421);
   U2084 : AO4 port map( A => n3557, B => n1147, C => n2450, D => n2341, Z => 
                           n5422);
   U2085 : AO4 port map( A => n3554, B => n1191, C => n365, D => n2340, Z => 
                           n5423);
   U2087 : AO4 port map( A => n3555, B => n1235, C => n365, D => n2339, Z => 
                           n5424);
   U2089 : AO4 port map( A => n3552, B => n442, C => n365, D => n2338, Z => 
                           n5425);
   U2091 : AO4 port map( A => n3553, B => n443, C => n365, D => n2337, Z => 
                           n5426);
   U2092 : AO4 port map( A => n3550, B => n487, C => n365, D => n2336, Z => 
                           n5427);
   U2094 : AO4 port map( A => n3551, B => n531, C => n365, D => n2335, Z => 
                           n5428);
   U2095 : AO4 port map( A => n3564, B => n1279, C => n365, D => n2334, Z => 
                           n5429);
   U2096 : AO4 port map( A => n3565, B => n1323, C => n365, D => n2333, Z => 
                           n5430);
   U2097 : AO4 port map( A => n3562, B => n1367, C => n365, D => n2332, Z => 
                           n5431);
   U2101 : AO4 port map( A => n3563, B => n1411, C => n365, D => n2331, Z => 
                           n5432);
   U2102 : AO4 port map( A => n3560, B => n575, C => n365, D => n2330, Z => 
                           n5433);
   U2103 : AO4 port map( A => n3561, B => n619, C => n365, D => n2329, Z => 
                           n5434);
   U2104 : AO4 port map( A => n3558, B => n663, C => n365, D => n2328, Z => 
                           n5435);
   U2106 : AO4 port map( A => n3559, B => n707, C => n365, D => n2327, Z => 
                           n5436);
   U2107 : AO4 port map( A => n3644, B => n390, C => n325, D => n2382, Z => 
                           n5893);
   U2110 : AO4 port map( A => n3645, B => n399, C => n2458, D => n2381, Z => 
                           n5894);
   U2111 : AO4 port map( A => n3642, B => n400, C => n325, D => n2380, Z => 
                           n5895);
   U2112 : AO4 port map( A => n3643, B => n401, C => n2458, D => n2379, Z => 
                           n5896);
   U2114 : AO4 port map( A => n3640, B => n402, C => n325, D => n2378, Z => 
                           n5897);
   U2115 : AO4 port map( A => n3641, B => n403, C => n2458, D => n2377, Z => 
                           n5898);
   U2116 : AO4 port map( A => n3638, B => n404, C => n325, D => n2376, Z => 
                           n5899);
   U2117 : AO4 port map( A => n3639, B => n405, C => n2458, D => n2375, Z => 
                           n5900);
   U2118 : AO4 port map( A => n3652, B => n406, C => n325, D => n2374, Z => 
                           n5901);
   U2119 : AO4 port map( A => n3653, B => n411, C => n2458, D => n2373, Z => 
                           n5902);
   U2122 : AO4 port map( A => n3650, B => n412, C => n2458, D => n2372, Z => 
                           n5903);
   U2123 : AO4 port map( A => n3651, B => n413, C => n2458, D => n2371, Z => 
                           n5904);
   U2124 : AO4 port map( A => n3648, B => n414, C => n2458, D => n2370, Z => 
                           n5905);
   U2127 : AO4 port map( A => n3649, B => n415, C => n2458, D => n2369, Z => 
                           n5906);
   U2128 : AO4 port map( A => n3646, B => n416, C => n325, D => n2368, Z => 
                           n5907);
   U2130 : AO4 port map( A => n3647, B => n417, C => n2458, D => n2367, Z => 
                           n5908);
   U2131 : AO4 port map( A => n3660, B => n418, C => n2458, D => n2366, Z => 
                           n5909);
   U2133 : AO4 port map( A => n3661, B => n423, C => n325, D => n2365, Z => 
                           n5910);
   U2134 : AO4 port map( A => n3658, B => n424, C => n2458, D => n2364, Z => 
                           n5911);
   U2135 : AO4 port map( A => n3659, B => n425, C => n2458, D => n2363, Z => 
                           n5912);
   U2136 : AO4 port map( A => n3656, B => n426, C => n325, D => n2362, Z => 
                           n5913);
   U2140 : AO4 port map( A => n3657, B => n427, C => n2458, D => n2361, Z => 
                           n5914);
   U2141 : AO4 port map( A => n3654, B => n428, C => n2458, D => n2360, Z => 
                           n5915);
   U2143 : AO4 port map( A => n3655, B => n429, C => n325, D => n2359, Z => 
                           n5916);
   U2147 : AO4 port map( A => n3604, B => n751, C => n2458, D => n2358, Z => 
                           n5917);
   U2148 : AO4 port map( A => n3605, B => n795, C => n2458, D => n2357, Z => 
                           n5918);
   U2149 : AO4 port map( A => n3602, B => n839, C => n325, D => n2356, Z => 
                           n5919);
   U2152 : AO4 port map( A => n3603, B => n883, C => n2458, D => n2355, Z => 
                           n5920);
   U2153 : AO4 port map( A => n3600, B => n430, C => n325, D => n2354, Z => 
                           n5921);
   U2154 : AO4 port map( A => n3601, B => n435, C => n325, D => n2353, Z => 
                           n5922);
   U2156 : AO4 port map( A => n3598, B => n436, C => n325, D => n2352, Z => 
                           n5923);
   U2157 : AO4 port map( A => n3599, B => n437, C => n325, D => n2351, Z => 
                           n5924);
   U2159 : AO4 port map( A => n3612, B => n927, C => n325, D => n2350, Z => 
                           n5925);
   U2161 : AO4 port map( A => n3613, B => n971, C => n325, D => n2349, Z => 
                           n5926);
   U2163 : AO4 port map( A => n3610, B => n1015, C => n325, D => n2348, Z => 
                           n5927);
   U2164 : AO4 port map( A => n3611, B => n1059, C => n325, D => n2347, Z => 
                           n5928);
   U2165 : AO4 port map( A => n3608, B => n438, C => n325, D => n2346, Z => 
                           n5929);
   U2166 : AO4 port map( A => n3609, B => n439, C => n325, D => n2345, Z => 
                           n5930);
   U2167 : AO4 port map( A => n3606, B => n440, C => n325, D => n2344, Z => 
                           n5931);
   U2169 : AO4 port map( A => n3607, B => n441, C => n325, D => n2343, Z => 
                           n5932);
   U2170 : AO4 port map( A => n3620, B => n1103, C => n325, D => n2342, Z => 
                           n5933);
   U2172 : AO4 port map( A => n3621, B => n1147, C => n325, D => n2341, Z => 
                           n5934);
   U2173 : AO4 port map( A => n3618, B => n1191, C => n325, D => n2340, Z => 
                           n5935);
   U2175 : AO4 port map( A => n3619, B => n1235, C => n325, D => n2339, Z => 
                           n5936);
   U2176 : AO4 port map( A => n3616, B => n442, C => n325, D => n2338, Z => 
                           n5937);
   U2178 : AO4 port map( A => n3617, B => n443, C => n325, D => n2337, Z => 
                           n5938);
   U2179 : AO4 port map( A => n3614, B => n487, C => n325, D => n2336, Z => 
                           n5939);
   U2182 : AO4 port map( A => n3615, B => n531, C => n2458, D => n2335, Z => 
                           n5940);
   U2184 : AO4 port map( A => n3628, B => n1279, C => n2458, D => n2334, Z => 
                           n5941);
   U2185 : AO4 port map( A => n3629, B => n1323, C => n2458, D => n2333, Z => 
                           n5942);
   U2186 : AO4 port map( A => n3626, B => n1367, C => n2458, D => n2332, Z => 
                           n5943);
   U2188 : AO4 port map( A => n3627, B => n1411, C => n2458, D => n2331, Z => 
                           n5944);
   U2190 : AO4 port map( A => n3624, B => n575, C => n2458, D => n2330, Z => 
                           n5945);
   U2191 : AO4 port map( A => n3625, B => n619, C => n2458, D => n2329, Z => 
                           n5946);
   U2193 : AO4 port map( A => n3622, B => n663, C => n2458, D => n2328, Z => 
                           n5947);
   U2194 : AO4 port map( A => n3623, B => n707, C => n2458, D => n2327, Z => 
                           n5948);
   U2195 : AO4 port map( A => n3708, B => n390, C => n314, D => n2382, Z => 
                           n6405);
   U2196 : AO4 port map( A => n3709, B => n399, C => n2466, D => n2381, Z => 
                           n6406);
   U2200 : AO4 port map( A => n3706, B => n400, C => n314, D => n2380, Z => 
                           n6407);
   U2202 : AO4 port map( A => n3707, B => n401, C => n2466, D => n2379, Z => 
                           n6408);
   U2203 : AO4 port map( A => n3704, B => n402, C => n314, D => n2378, Z => 
                           n6409);
   U2206 : AO4 port map( A => n3705, B => n403, C => n2466, D => n2377, Z => 
                           n6410);
   U2207 : AO4 port map( A => n3702, B => n404, C => n314, D => n2376, Z => 
                           n6411);
   U2209 : AO4 port map( A => n3703, B => n405, C => n2466, D => n2375, Z => 
                           n6412);
   U2211 : AO4 port map( A => n3716, B => n406, C => n314, D => n2374, Z => 
                           n6413);
   U2217 : AO4 port map( A => n3717, B => n411, C => n2466, D => n2373, Z => 
                           n6414);
   U2218 : AO4 port map( A => n3714, B => n412, C => n2466, D => n2372, Z => 
                           n6415);
   U2219 : AO4 port map( A => n3715, B => n413, C => n2466, D => n2371, Z => 
                           n6416);
   U2220 : AO4 port map( A => n3712, B => n414, C => n2466, D => n2370, Z => 
                           n6417);
   U2221 : AO4 port map( A => n3713, B => n415, C => n2466, D => n2369, Z => 
                           n6418);
   U2225 : AO4 port map( A => n3710, B => n416, C => n314, D => n2368, Z => 
                           n6419);
   U2226 : AO4 port map( A => n3711, B => n417, C => n2466, D => n2367, Z => 
                           n6420);
   U2228 : AO4 port map( A => n3724, B => n418, C => n2466, D => n2366, Z => 
                           n6421);
   U2230 : AO4 port map( A => n3725, B => n423, C => n314, D => n2365, Z => 
                           n6422);
   U2232 : AO4 port map( A => n3722, B => n424, C => n2466, D => n2364, Z => 
                           n6423);
   U2233 : AO4 port map( A => n3723, B => n425, C => n2466, D => n2363, Z => 
                           n6424);
   U2236 : AO4 port map( A => n3720, B => n426, C => n314, D => n2362, Z => 
                           n6425);
   U2241 : AO4 port map( A => n3721, B => n427, C => n2466, D => n2361, Z => 
                           n6426);
   U2242 : AO4 port map( A => n3718, B => n428, C => n2466, D => n2360, Z => 
                           n6427);
   U2244 : AO4 port map( A => n3719, B => n429, C => n314, D => n2359, Z => 
                           n6428);
   U2246 : AO4 port map( A => n3668, B => n751, C => n2466, D => n2358, Z => 
                           n6429);
   U2247 : AO4 port map( A => n3669, B => n795, C => n2466, D => n2357, Z => 
                           n6430);
   U2248 : AO4 port map( A => n3666, B => n839, C => n314, D => n2356, Z => 
                           n6431);
   U2251 : AO4 port map( A => n3667, B => n883, C => n2466, D => n2355, Z => 
                           n6432);
   U2252 : AO4 port map( A => n3664, B => n430, C => n314, D => n2354, Z => 
                           n6433);
   U2257 : AO4 port map( A => n3665, B => n435, C => n314, D => n2353, Z => 
                           n6434);
   U2259 : AO4 port map( A => n3662, B => n436, C => n314, D => n2352, Z => 
                           n6435);
   U2260 : AO4 port map( A => n3663, B => n437, C => n314, D => n2351, Z => 
                           n6436);
   U2262 : AO4 port map( A => n3676, B => n927, C => n314, D => n2350, Z => 
                           n6437);
   U2267 : AO4 port map( A => n3677, B => n971, C => n314, D => n2349, Z => 
                           n6438);
   U2269 : AO4 port map( A => n3674, B => n1015, C => n314, D => n2348, Z => 
                           n6439);
   U2272 : AO4 port map( A => n3675, B => n1059, C => n314, D => n2347, Z => 
                           n6440);
   U2275 : AO4 port map( A => n3672, B => n438, C => n314, D => n2346, Z => 
                           n6441);
   U2277 : AO4 port map( A => n3673, B => n439, C => n314, D => n2345, Z => 
                           n6442);
   U2278 : AO4 port map( A => n3670, B => n440, C => n314, D => n2344, Z => 
                           n6443);
   U2283 : AO4 port map( A => n3671, B => n441, C => n314, D => n2343, Z => 
                           n6444);
   U2285 : AO4 port map( A => n3684, B => n1103, C => n314, D => n2342, Z => 
                           n6445);
   U2288 : AO4 port map( A => n3685, B => n1147, C => n314, D => n2341, Z => 
                           n6446);
   U2291 : AO4 port map( A => n3682, B => n1191, C => n314, D => n2340, Z => 
                           n6447);
   U2293 : AO4 port map( A => n3683, B => n1235, C => n314, D => n2339, Z => 
                           n6448);
   U2296 : AO4 port map( A => n3680, B => n442, C => n314, D => n2338, Z => 
                           n6449);
   U2300 : AO4 port map( A => n3681, B => n443, C => n314, D => n2337, Z => 
                           n6450);
   U2301 : AO4 port map( A => n3678, B => n487, C => n314, D => n2336, Z => 
                           n6451);
   U2302 : AO4 port map( A => n3679, B => n531, C => n2466, D => n2335, Z => 
                           n6452);
   U2304 : AO4 port map( A => n3692, B => n1279, C => n2466, D => n2334, Z => 
                           n6453);
   U2307 : AO4 port map( A => n3693, B => n1323, C => n2466, D => n2333, Z => 
                           n6454);
   U2308 : AO4 port map( A => n3690, B => n1367, C => n2466, D => n2332, Z => 
                           n6455);
   U2310 : AO4 port map( A => n3691, B => n1411, C => n2466, D => n2331, Z => 
                           n6456);
   U2312 : AO4 port map( A => n3688, B => n575, C => n2466, D => n2330, Z => 
                           n6457);
   U2313 : AO4 port map( A => n3689, B => n619, C => n2466, D => n2329, Z => 
                           n6458);
   U2315 : AO4 port map( A => n3686, B => n663, C => n2466, D => n2328, Z => 
                           n6459);
   U2317 : AO4 port map( A => n3687, B => n707, C => n2466, D => n2327, Z => 
                           n6460);
   U2318 : AO4 port map( A => n3772, B => n390, C => n364, D => n2382, Z => 
                           n4869);
   U2319 : AO4 port map( A => n3773, B => n399, C => n2442, D => n2381, Z => 
                           n4870);
   U2321 : AO4 port map( A => n3770, B => n400, C => n364, D => n2380, Z => 
                           n4871);
   U2322 : AO4 port map( A => n3771, B => n401, C => n2442, D => n2379, Z => 
                           n4872);
   U2323 : AO4 port map( A => n3768, B => n402, C => n364, D => n2378, Z => 
                           n4873);
   U2324 : AO4 port map( A => n3769, B => n403, C => n2442, D => n2377, Z => 
                           n4874);
   U2326 : AO4 port map( A => n3766, B => n404, C => n364, D => n2376, Z => 
                           n4875);
   U2327 : AO4 port map( A => n3767, B => n405, C => n2442, D => n2375, Z => 
                           n4876);
   U2330 : AO4 port map( A => n3780, B => n406, C => n364, D => n2374, Z => 
                           n4877);
   U2332 : AO4 port map( A => n3781, B => n411, C => n2442, D => n2373, Z => 
                           n4878);
   U2334 : AO4 port map( A => n3778, B => n412, C => n2442, D => n2372, Z => 
                           n4879);
   U2335 : AO4 port map( A => n3779, B => n413, C => n2442, D => n2371, Z => 
                           n4880);
   U2336 : AO4 port map( A => n3776, B => n414, C => n2442, D => n2370, Z => 
                           n4881);
   U2338 : AO4 port map( A => n3777, B => n415, C => n2442, D => n2369, Z => 
                           n4882);
   U2340 : AO4 port map( A => n3774, B => n416, C => n364, D => n2368, Z => 
                           n4883);
   U2341 : AO4 port map( A => n3775, B => n417, C => n2442, D => n2367, Z => 
                           n4884);
   U2342 : AO4 port map( A => n3788, B => n418, C => n2442, D => n2366, Z => 
                           n4885);
   U2343 : AO4 port map( A => n3789, B => n423, C => n364, D => n2365, Z => 
                           n4886);
   U2344 : AO4 port map( A => n3786, B => n424, C => n2442, D => n2364, Z => 
                           n4887);
   U2345 : AO4 port map( A => n3787, B => n425, C => n2442, D => n2363, Z => 
                           n4888);
   U2348 : AO4 port map( A => n3784, B => n426, C => n364, D => n2362, Z => 
                           n4889);
   U2349 : AO4 port map( A => n3785, B => n427, C => n2442, D => n2361, Z => 
                           n4890);
   U2351 : AO4 port map( A => n3782, B => n428, C => n2442, D => n2360, Z => 
                           n4891);
   U2352 : AO4 port map( A => n3783, B => n429, C => n364, D => n2359, Z => 
                           n4892);
   U2354 : AO4 port map( A => n3732, B => n751, C => n2442, D => n2358, Z => 
                           n4893);
   U2356 : AO4 port map( A => n3733, B => n795, C => n2442, D => n2357, Z => 
                           n4894);
   U2357 : AO4 port map( A => n3730, B => n839, C => n364, D => n2356, Z => 
                           n4895);
   U2359 : AO4 port map( A => n3731, B => n883, C => n2442, D => n2355, Z => 
                           n4896);
   U2360 : AO4 port map( A => n3728, B => n430, C => n364, D => n2354, Z => 
                           n4897);
   U2365 : AO4 port map( A => n3729, B => n435, C => n364, D => n2353, Z => 
                           n4898);
   U2366 : AO4 port map( A => n3726, B => n436, C => n364, D => n2352, Z => 
                           n4899);
   U2367 : AO4 port map( A => n3727, B => n437, C => n364, D => n2351, Z => 
                           n4900);
   U2368 : AO4 port map( A => n3740, B => n927, C => n364, D => n2350, Z => 
                           n4901);
   U2369 : AO4 port map( A => n3741, B => n971, C => n364, D => n2349, Z => 
                           n4902);
   U2371 : AO4 port map( A => n3738, B => n1015, C => n364, D => n2348, Z => 
                           n4903);
   U2372 : AO4 port map( A => n3739, B => n1059, C => n364, D => n2347, Z => 
                           n4904);
   U2373 : AO4 port map( A => n3736, B => n438, C => n364, D => n2346, Z => 
                           n4905);
   U2374 : AO4 port map( A => n3737, B => n439, C => n364, D => n2345, Z => 
                           n4906);
   U2375 : AO4 port map( A => n3734, B => n440, C => n364, D => n2344, Z => 
                           n4907);
   U2376 : AO4 port map( A => n3735, B => n441, C => n364, D => n2343, Z => 
                           n4908);
   U2377 : AO4 port map( A => n3748, B => n1103, C => n364, D => n2342, Z => 
                           n4909);
   U2378 : AO4 port map( A => n3749, B => n1147, C => n364, D => n2341, Z => 
                           n4910);
   U2379 : AO4 port map( A => n3746, B => n1191, C => n364, D => n2340, Z => 
                           n4911);
   U2380 : AO4 port map( A => n3747, B => n1235, C => n364, D => n2339, Z => 
                           n4912);
   U2381 : AO4 port map( A => n3744, B => n442, C => n364, D => n2338, Z => 
                           n4913);
   U2382 : AO4 port map( A => n3745, B => n443, C => n364, D => n2337, Z => 
                           n4914);
   U2383 : AO4 port map( A => n3742, B => n487, C => n364, D => n2336, Z => 
                           n4915);
   U2384 : AO4 port map( A => n3743, B => n531, C => n2442, D => n2335, Z => 
                           n4916);
   U2385 : AO4 port map( A => n3756, B => n1279, C => n2442, D => n2334, Z => 
                           n4917);
   U2386 : AO4 port map( A => n3757, B => n1323, C => n2442, D => n2333, Z => 
                           n4918);
   U2387 : AO4 port map( A => n3754, B => n1367, C => n2442, D => n2332, Z => 
                           n4919);
   U2388 : AO4 port map( A => n3755, B => n1411, C => n2442, D => n2331, Z => 
                           n4920);
   U2389 : AO4 port map( A => n3752, B => n575, C => n2442, D => n2330, Z => 
                           n4921);
   U2390 : AO4 port map( A => n3753, B => n619, C => n2442, D => n2329, Z => 
                           n4922);
   U2391 : AO4 port map( A => n3750, B => n663, C => n2442, D => n2328, Z => 
                           n4923);
   U2392 : AO4 port map( A => n3751, B => n707, C => n2442, D => n2327, Z => 
                           n4924);
   U2393 : AO4 port map( A => n3836, B => n390, C => n363, D => n2382, Z => 
                           n5445);
   U2394 : AO4 port map( A => n3837, B => n399, C => n2451, D => n2381, Z => 
                           n5446);
   U2395 : AO4 port map( A => n3834, B => n400, C => n363, D => n2380, Z => 
                           n5447);
   U2396 : AO4 port map( A => n3835, B => n401, C => n2451, D => n2379, Z => 
                           n5448);
   U2397 : AO4 port map( A => n3832, B => n402, C => n363, D => n2378, Z => 
                           n5449);
   U2398 : AO4 port map( A => n3833, B => n403, C => n2451, D => n2377, Z => 
                           n5450);
   U2399 : AO4 port map( A => n3830, B => n404, C => n363, D => n2376, Z => 
                           n5451);
   U2400 : AO4 port map( A => n3831, B => n405, C => n2451, D => n2375, Z => 
                           n5452);
   U2401 : AO4 port map( A => n3844, B => n406, C => n363, D => n2374, Z => 
                           n5453);
   U2402 : AO4 port map( A => n3845, B => n411, C => n2451, D => n2373, Z => 
                           n5454);
   U2403 : AO4 port map( A => n3842, B => n412, C => n2451, D => n2372, Z => 
                           n5455);
   U2404 : AO4 port map( A => n3843, B => n413, C => n2451, D => n2371, Z => 
                           n5456);
   U2405 : AO4 port map( A => n3840, B => n414, C => n2451, D => n2370, Z => 
                           n5457);
   U2406 : AO4 port map( A => n3841, B => n415, C => n2451, D => n2369, Z => 
                           n5458);
   U2407 : AO4 port map( A => n3838, B => n416, C => n363, D => n2368, Z => 
                           n5459);
   U2408 : AO4 port map( A => n3839, B => n417, C => n2451, D => n2367, Z => 
                           n5460);
   U2409 : AO4 port map( A => n3852, B => n418, C => n2451, D => n2366, Z => 
                           n5461);
   U2410 : AO4 port map( A => n3853, B => n423, C => n363, D => n2365, Z => 
                           n5462);
   U2411 : AO4 port map( A => n3850, B => n424, C => n2451, D => n2364, Z => 
                           n5463);
   U2412 : AO4 port map( A => n3851, B => n425, C => n2451, D => n2363, Z => 
                           n5464);
   U2413 : AO4 port map( A => n3848, B => n426, C => n363, D => n2362, Z => 
                           n5465);
   U2414 : AO4 port map( A => n3849, B => n427, C => n2451, D => n2361, Z => 
                           n5466);
   U2415 : AO4 port map( A => n3846, B => n428, C => n2451, D => n2360, Z => 
                           n5467);
   U2416 : AO4 port map( A => n3847, B => n429, C => n363, D => n2359, Z => 
                           n5468);
   U2417 : AO4 port map( A => n3796, B => n751, C => n2451, D => n2358, Z => 
                           n5469);
   U2418 : AO4 port map( A => n3797, B => n795, C => n2451, D => n2357, Z => 
                           n5470);
   U2419 : AO4 port map( A => n3794, B => n839, C => n363, D => n2356, Z => 
                           n5471);
   U2420 : AO4 port map( A => n3795, B => n883, C => n2451, D => n2355, Z => 
                           n5472);
   U2421 : AO4 port map( A => n3792, B => n430, C => n363, D => n2354, Z => 
                           n5473);
   U2422 : AO4 port map( A => n3793, B => n435, C => n363, D => n2353, Z => 
                           n5474);
   U2423 : AO4 port map( A => n3790, B => n436, C => n363, D => n2352, Z => 
                           n5475);
   U2424 : AO4 port map( A => n3791, B => n437, C => n363, D => n2351, Z => 
                           n5476);
   U2425 : AO4 port map( A => n3804, B => n927, C => n363, D => n2350, Z => 
                           n5477);
   U2426 : AO4 port map( A => n3805, B => n971, C => n363, D => n2349, Z => 
                           n5478);
   U2427 : AO4 port map( A => n3802, B => n1015, C => n363, D => n2348, Z => 
                           n5479);
   U2428 : AO4 port map( A => n3803, B => n1059, C => n363, D => n2347, Z => 
                           n5480);
   U2429 : AO4 port map( A => n3800, B => n438, C => n363, D => n2346, Z => 
                           n5481);
   U2430 : AO4 port map( A => n3801, B => n439, C => n363, D => n2345, Z => 
                           n5482);
   U2431 : AO4 port map( A => n3798, B => n440, C => n363, D => n2344, Z => 
                           n5483);
   U2432 : AO4 port map( A => n3799, B => n441, C => n363, D => n2343, Z => 
                           n5484);
   U2433 : AO4 port map( A => n3812, B => n1103, C => n363, D => n2342, Z => 
                           n5485);
   U2434 : AO4 port map( A => n3813, B => n1147, C => n363, D => n2341, Z => 
                           n5486);
   U2435 : AO4 port map( A => n3810, B => n1191, C => n363, D => n2340, Z => 
                           n5487);
   U2436 : AO4 port map( A => n3811, B => n1235, C => n363, D => n2339, Z => 
                           n5488);
   U2437 : AO4 port map( A => n3808, B => n442, C => n363, D => n2338, Z => 
                           n5489);
   U2438 : AO4 port map( A => n3809, B => n443, C => n363, D => n2337, Z => 
                           n5490);
   U2439 : AO4 port map( A => n3806, B => n487, C => n363, D => n2336, Z => 
                           n5491);
   U2440 : AO4 port map( A => n3807, B => n531, C => n2451, D => n2335, Z => 
                           n5492);
   U2441 : AO4 port map( A => n3820, B => n1279, C => n2451, D => n2334, Z => 
                           n5493);
   U2442 : AO4 port map( A => n3821, B => n1323, C => n2451, D => n2333, Z => 
                           n5494);
   U2443 : AO4 port map( A => n3818, B => n1367, C => n2451, D => n2332, Z => 
                           n5495);
   U2444 : AO4 port map( A => n3819, B => n1411, C => n2451, D => n2331, Z => 
                           n5496);
   U2445 : AO4 port map( A => n3816, B => n575, C => n2451, D => n2330, Z => 
                           n5497);
   U2446 : AO4 port map( A => n3817, B => n619, C => n2451, D => n2329, Z => 
                           n5498);
   U2447 : AO4 port map( A => n3814, B => n663, C => n2451, D => n2328, Z => 
                           n5499);
   U2448 : AO4 port map( A => n3815, B => n707, C => n2451, D => n2327, Z => 
                           n5500);
   U2449 : AO4 port map( A => n3900, B => n390, C => n2459, D => n2382, Z => 
                           n5957);
   U2450 : AO4 port map( A => n3901, B => n399, C => n2459, D => n2381, Z => 
                           n5958);
   U2451 : AO4 port map( A => n3898, B => n400, C => n2459, D => n2380, Z => 
                           n5959);
   U2452 : AO4 port map( A => n3899, B => n401, C => n2459, D => n2379, Z => 
                           n5960);
   U2453 : AO4 port map( A => n3896, B => n402, C => n2459, D => n2378, Z => 
                           n5961);
   U2454 : AO4 port map( A => n3897, B => n403, C => n2459, D => n2377, Z => 
                           n5962);
   U2455 : AO4 port map( A => n3894, B => n404, C => n2459, D => n2376, Z => 
                           n5963);
   U2456 : AO4 port map( A => n3895, B => n405, C => n2459, D => n2375, Z => 
                           n5964);
   U2457 : AO4 port map( A => n3908, B => n406, C => n303, D => n2374, Z => 
                           n5965);
   U2458 : AO4 port map( A => n3909, B => n411, C => n2459, D => n2373, Z => 
                           n5966);
   U2459 : AO4 port map( A => n3906, B => n412, C => n2459, D => n2372, Z => 
                           n5967);
   U2460 : AO4 port map( A => n3907, B => n413, C => n2459, D => n2371, Z => 
                           n5968);
   U2461 : AO4 port map( A => n3904, B => n414, C => n303, D => n2370, Z => 
                           n5969);
   U2462 : AO4 port map( A => n3905, B => n415, C => n2459, D => n2369, Z => 
                           n5970);
   U2463 : AO4 port map( A => n3902, B => n416, C => n303, D => n2368, Z => 
                           n5971);
   U2464 : AO4 port map( A => n3903, B => n417, C => n303, D => n2367, Z => 
                           n5972);
   U2465 : AO4 port map( A => n3916, B => n418, C => n303, D => n2366, Z => 
                           n5973);
   U2466 : AO4 port map( A => n3917, B => n423, C => n303, D => n2365, Z => 
                           n5974);
   U2467 : AO4 port map( A => n3914, B => n424, C => n303, D => n2364, Z => 
                           n5975);
   U2468 : AO4 port map( A => n3915, B => n425, C => n303, D => n2363, Z => 
                           n5976);
   U2469 : AO4 port map( A => n3912, B => n426, C => n303, D => n2362, Z => 
                           n5977);
   U2470 : AO4 port map( A => n3913, B => n427, C => n303, D => n2361, Z => 
                           n5978);
   U2471 : AO4 port map( A => n3910, B => n428, C => n303, D => n2360, Z => 
                           n5979);
   U2472 : AO4 port map( A => n3911, B => n429, C => n303, D => n2359, Z => 
                           n5980);
   U2473 : AO4 port map( A => n3860, B => n751, C => n303, D => n2358, Z => 
                           n5981);
   U2474 : AO4 port map( A => n3861, B => n795, C => n303, D => n2357, Z => 
                           n5982);
   U2475 : AO4 port map( A => n3858, B => n839, C => n303, D => n2356, Z => 
                           n5983);
   U2476 : AO4 port map( A => n3859, B => n883, C => n303, D => n2355, Z => 
                           n5984);
   U2477 : AO4 port map( A => n3856, B => n430, C => n303, D => n2354, Z => 
                           n5985);
   U2478 : AO4 port map( A => n3857, B => n435, C => n303, D => n2353, Z => 
                           n5986);
   U2479 : AO4 port map( A => n3854, B => n436, C => n303, D => n2352, Z => 
                           n5987);
   U2480 : AO4 port map( A => n3855, B => n437, C => n303, D => n2351, Z => 
                           n5988);
   U2481 : AO4 port map( A => n3868, B => n927, C => n303, D => n2350, Z => 
                           n5989);
   U2482 : AO4 port map( A => n3869, B => n971, C => n303, D => n2349, Z => 
                           n5990);
   U2483 : AO4 port map( A => n3866, B => n1015, C => n303, D => n2348, Z => 
                           n5991);
   U2484 : AO4 port map( A => n3867, B => n1059, C => n303, D => n2347, Z => 
                           n5992);
   U2485 : AO4 port map( A => n3864, B => n438, C => n303, D => n2346, Z => 
                           n5993);
   U2486 : AO4 port map( A => n3865, B => n439, C => n303, D => n2345, Z => 
                           n5994);
   U2487 : AO4 port map( A => n3862, B => n440, C => n2459, D => n2344, Z => 
                           n5995);
   U2488 : AO4 port map( A => n3863, B => n441, C => n2459, D => n2343, Z => 
                           n5996);
   U2489 : AO4 port map( A => n3876, B => n1103, C => n2459, D => n2342, Z => 
                           n5997);
   U2490 : AO4 port map( A => n3877, B => n1147, C => n2459, D => n2341, Z => 
                           n5998);
   U2491 : AO4 port map( A => n3874, B => n1191, C => n2459, D => n2340, Z => 
                           n5999);
   U2492 : AO4 port map( A => n3875, B => n1235, C => n303, D => n2339, Z => 
                           n6000);
   U2493 : AO4 port map( A => n3872, B => n442, C => n2459, D => n2338, Z => 
                           n6001);
   U2494 : AO4 port map( A => n3873, B => n443, C => n2459, D => n2337, Z => 
                           n6002);
   U2495 : AO4 port map( A => n3870, B => n487, C => n303, D => n2336, Z => 
                           n6003);
   U2496 : AO4 port map( A => n3871, B => n531, C => n2459, D => n2335, Z => 
                           n6004);
   U2497 : AO4 port map( A => n3884, B => n1279, C => n2459, D => n2334, Z => 
                           n6005);
   U2498 : AO4 port map( A => n3885, B => n1323, C => n303, D => n2333, Z => 
                           n6006);
   U2499 : AO4 port map( A => n3882, B => n1367, C => n2459, D => n2332, Z => 
                           n6007);
   U2500 : AO4 port map( A => n3883, B => n1411, C => n2459, D => n2331, Z => 
                           n6008);
   U2501 : AO4 port map( A => n3880, B => n575, C => n303, D => n2330, Z => 
                           n6009);
   U2502 : AO4 port map( A => n3881, B => n619, C => n2459, D => n2329, Z => 
                           n6010);
   U2503 : AO4 port map( A => n3878, B => n663, C => n2459, D => n2328, Z => 
                           n6011);
   U2504 : AO4 port map( A => n3879, B => n707, C => n303, D => n2327, Z => 
                           n6012);
   U2505 : AO4 port map( A => n3964, B => n390, C => n301, D => n2382, Z => 
                           n6469);
   U2506 : AO4 port map( A => n3965, B => n399, C => n2467, D => n2381, Z => 
                           n6470);
   U2507 : AO4 port map( A => n3962, B => n400, C => n301, D => n2380, Z => 
                           n6471);
   U2508 : AO4 port map( A => n3963, B => n401, C => n2467, D => n2379, Z => 
                           n6472);
   U2509 : AO4 port map( A => n3960, B => n402, C => n301, D => n2378, Z => 
                           n6473);
   U2510 : AO4 port map( A => n3961, B => n403, C => n2467, D => n2377, Z => 
                           n6474);
   U2511 : AO4 port map( A => n3958, B => n404, C => n301, D => n2376, Z => 
                           n6475);
   U2512 : AO4 port map( A => n3959, B => n405, C => n2467, D => n2375, Z => 
                           n6476);
   U2513 : AO4 port map( A => n3972, B => n406, C => n301, D => n2374, Z => 
                           n6477);
   U2514 : AO4 port map( A => n3973, B => n411, C => n2467, D => n2373, Z => 
                           n6478);
   U2515 : AO4 port map( A => n3970, B => n412, C => n2467, D => n2372, Z => 
                           n6479);
   U2516 : AO4 port map( A => n3971, B => n413, C => n2467, D => n2371, Z => 
                           n6480);
   U2517 : AO4 port map( A => n3968, B => n414, C => n2467, D => n2370, Z => 
                           n6481);
   U2518 : AO4 port map( A => n3969, B => n415, C => n2467, D => n2369, Z => 
                           n6482);
   U2519 : AO4 port map( A => n3966, B => n416, C => n301, D => n2368, Z => 
                           n6483);
   U2520 : AO4 port map( A => n3967, B => n417, C => n2467, D => n2367, Z => 
                           n6484);
   U2521 : AO4 port map( A => n3980, B => n418, C => n2467, D => n2366, Z => 
                           n6485);
   U2522 : AO4 port map( A => n3981, B => n423, C => n301, D => n2365, Z => 
                           n6486);
   U2523 : AO4 port map( A => n3978, B => n424, C => n2467, D => n2364, Z => 
                           n6487);
   U2524 : AO4 port map( A => n3979, B => n425, C => n2467, D => n2363, Z => 
                           n6488);
   U2525 : AO4 port map( A => n3976, B => n426, C => n301, D => n2362, Z => 
                           n6489);
   U2526 : AO4 port map( A => n3977, B => n427, C => n2467, D => n2361, Z => 
                           n6490);
   U2527 : AO4 port map( A => n3974, B => n428, C => n2467, D => n2360, Z => 
                           n6491);
   U2528 : AO4 port map( A => n3975, B => n429, C => n301, D => n2359, Z => 
                           n6492);
   U2529 : AO4 port map( A => n3924, B => n751, C => n2467, D => n2358, Z => 
                           n6493);
   U2530 : AO4 port map( A => n3925, B => n795, C => n2467, D => n2357, Z => 
                           n6494);
   U2531 : AO4 port map( A => n3922, B => n839, C => n301, D => n2356, Z => 
                           n6495);
   U2532 : AO4 port map( A => n3923, B => n883, C => n2467, D => n2355, Z => 
                           n6496);
   U2533 : AO4 port map( A => n3920, B => n430, C => n301, D => n2354, Z => 
                           n6497);
   U2534 : AO4 port map( A => n3921, B => n435, C => n301, D => n2353, Z => 
                           n6498);
   U2535 : AO4 port map( A => n3918, B => n436, C => n301, D => n2352, Z => 
                           n6499);
   U2536 : AO4 port map( A => n3919, B => n437, C => n301, D => n2351, Z => 
                           n6500);
   U2537 : AO4 port map( A => n3932, B => n927, C => n301, D => n2350, Z => 
                           n6501);
   U2538 : AO4 port map( A => n3933, B => n971, C => n301, D => n2349, Z => 
                           n6502);
   U2539 : AO4 port map( A => n3930, B => n1015, C => n301, D => n2348, Z => 
                           n6503);
   U2540 : AO4 port map( A => n3931, B => n1059, C => n301, D => n2347, Z => 
                           n6504);
   U2541 : AO4 port map( A => n3928, B => n438, C => n301, D => n2346, Z => 
                           n6505);
   U2542 : AO4 port map( A => n3929, B => n439, C => n301, D => n2345, Z => 
                           n6506);
   U2543 : AO4 port map( A => n3926, B => n440, C => n301, D => n2344, Z => 
                           n6507);
   U2544 : AO4 port map( A => n3927, B => n441, C => n301, D => n2343, Z => 
                           n6508);
   U2545 : AO4 port map( A => n3940, B => n1103, C => n301, D => n2342, Z => 
                           n6509);
   U2546 : AO4 port map( A => n3941, B => n1147, C => n301, D => n2341, Z => 
                           n6510);
   U2547 : AO4 port map( A => n3938, B => n1191, C => n301, D => n2340, Z => 
                           n6511);
   U2548 : AO4 port map( A => n3939, B => n1235, C => n301, D => n2339, Z => 
                           n6512);
   U2549 : AO4 port map( A => n3936, B => n442, C => n301, D => n2338, Z => 
                           n6513);
   U2550 : AO4 port map( A => n3937, B => n443, C => n301, D => n2337, Z => 
                           n6514);
   U2551 : AO4 port map( A => n3934, B => n487, C => n301, D => n2336, Z => 
                           n6515);
   U2552 : AO4 port map( A => n3935, B => n531, C => n2467, D => n2335, Z => 
                           n6516);
   U2553 : AO4 port map( A => n3948, B => n1279, C => n2467, D => n2334, Z => 
                           n6517);
   U2554 : AO4 port map( A => n3949, B => n1323, C => n2467, D => n2333, Z => 
                           n6518);
   U2555 : AO4 port map( A => n3946, B => n1367, C => n2467, D => n2332, Z => 
                           n6519);
   U2556 : AO4 port map( A => n3947, B => n1411, C => n2467, D => n2331, Z => 
                           n6520);
   U2557 : AO4 port map( A => n3944, B => n575, C => n2467, D => n2330, Z => 
                           n6521);
   U2558 : AO4 port map( A => n3945, B => n619, C => n2467, D => n2329, Z => 
                           n6522);
   U2559 : AO4 port map( A => n3942, B => n663, C => n2467, D => n2328, Z => 
                           n6523);
   U2560 : AO4 port map( A => n3943, B => n707, C => n2467, D => n2327, Z => 
                           n6524);
   U2561 : AO4 port map( A => n4028, B => n390, C => n2443, D => n2382, Z => 
                           n4933);
   U2562 : AO4 port map( A => n4029, B => n399, C => n2443, D => n2381, Z => 
                           n4934);
   U2563 : AO4 port map( A => n4026, B => n400, C => n2443, D => n2380, Z => 
                           n4935);
   U2564 : AO4 port map( A => n4027, B => n401, C => n2443, D => n2379, Z => 
                           n4936);
   U2565 : AO4 port map( A => n4024, B => n402, C => n2443, D => n2378, Z => 
                           n4937);
   U2566 : AO4 port map( A => n4025, B => n403, C => n2443, D => n2377, Z => 
                           n4938);
   U2567 : AO4 port map( A => n4022, B => n404, C => n2443, D => n2376, Z => 
                           n4939);
   U2568 : AO4 port map( A => n4023, B => n405, C => n2443, D => n2375, Z => 
                           n4940);
   U2569 : AO4 port map( A => n4036, B => n406, C => n362, D => n2374, Z => 
                           n4941);
   U2570 : AO4 port map( A => n4037, B => n411, C => n2443, D => n2373, Z => 
                           n4942);
   U2571 : AO4 port map( A => n4034, B => n412, C => n2443, D => n2372, Z => 
                           n4943);
   U2572 : AO4 port map( A => n4035, B => n413, C => n2443, D => n2371, Z => 
                           n4944);
   U2573 : AO4 port map( A => n4032, B => n414, C => n362, D => n2370, Z => 
                           n4945);
   U2574 : AO4 port map( A => n4033, B => n415, C => n2443, D => n2369, Z => 
                           n4946);
   U2575 : AO4 port map( A => n4030, B => n416, C => n362, D => n2368, Z => 
                           n4947);
   U2576 : AO4 port map( A => n4031, B => n417, C => n362, D => n2367, Z => 
                           n4948);
   U2577 : AO4 port map( A => n4044, B => n418, C => n362, D => n2366, Z => 
                           n4949);
   U2578 : AO4 port map( A => n4045, B => n423, C => n362, D => n2365, Z => 
                           n4950);
   U2579 : AO4 port map( A => n4042, B => n424, C => n362, D => n2364, Z => 
                           n4951);
   U2580 : AO4 port map( A => n4043, B => n425, C => n362, D => n2363, Z => 
                           n4952);
   U2581 : AO4 port map( A => n4040, B => n426, C => n362, D => n2362, Z => 
                           n4953);
   U2582 : AO4 port map( A => n4041, B => n427, C => n362, D => n2361, Z => 
                           n4954);
   U2583 : AO4 port map( A => n4038, B => n428, C => n362, D => n2360, Z => 
                           n4955);
   U2584 : AO4 port map( A => n4039, B => n429, C => n362, D => n2359, Z => 
                           n4956);
   U2585 : AO4 port map( A => n3988, B => n751, C => n362, D => n2358, Z => 
                           n4957);
   U2586 : AO4 port map( A => n3989, B => n795, C => n362, D => n2357, Z => 
                           n4958);
   U2587 : AO4 port map( A => n3986, B => n839, C => n362, D => n2356, Z => 
                           n4959);
   U2588 : AO4 port map( A => n3987, B => n883, C => n362, D => n2355, Z => 
                           n4960);
   U2589 : AO4 port map( A => n3984, B => n430, C => n362, D => n2354, Z => 
                           n4961);
   U2590 : AO4 port map( A => n3985, B => n435, C => n362, D => n2353, Z => 
                           n4962);
   U2591 : AO4 port map( A => n3982, B => n436, C => n362, D => n2352, Z => 
                           n4963);
   U2592 : AO4 port map( A => n3983, B => n437, C => n362, D => n2351, Z => 
                           n4964);
   U2593 : AO4 port map( A => n3996, B => n927, C => n362, D => n2350, Z => 
                           n4965);
   U2594 : AO4 port map( A => n3997, B => n971, C => n362, D => n2349, Z => 
                           n4966);
   U2595 : AO4 port map( A => n3994, B => n1015, C => n362, D => n2348, Z => 
                           n4967);
   U2596 : AO4 port map( A => n3995, B => n1059, C => n362, D => n2347, Z => 
                           n4968);
   U2597 : AO4 port map( A => n3992, B => n438, C => n362, D => n2346, Z => 
                           n4969);
   U2598 : AO4 port map( A => n3993, B => n439, C => n362, D => n2345, Z => 
                           n4970);
   U2599 : AO4 port map( A => n3990, B => n440, C => n2443, D => n2344, Z => 
                           n4971);
   U2600 : AO4 port map( A => n3991, B => n441, C => n2443, D => n2343, Z => 
                           n4972);
   U2601 : AO4 port map( A => n4004, B => n1103, C => n2443, D => n2342, Z => 
                           n4973);
   U2602 : AO4 port map( A => n4005, B => n1147, C => n2443, D => n2341, Z => 
                           n4974);
   U2603 : AO4 port map( A => n4002, B => n1191, C => n2443, D => n2340, Z => 
                           n4975);
   U2604 : AO4 port map( A => n4003, B => n1235, C => n362, D => n2339, Z => 
                           n4976);
   U2605 : AO4 port map( A => n4000, B => n442, C => n2443, D => n2338, Z => 
                           n4977);
   U2606 : AO4 port map( A => n4001, B => n443, C => n2443, D => n2337, Z => 
                           n4978);
   U2607 : AO4 port map( A => n3998, B => n487, C => n362, D => n2336, Z => 
                           n4979);
   U2608 : AO4 port map( A => n3999, B => n531, C => n2443, D => n2335, Z => 
                           n4980);
   U2609 : AO4 port map( A => n4012, B => n1279, C => n2443, D => n2334, Z => 
                           n4981);
   U2610 : AO4 port map( A => n4013, B => n1323, C => n362, D => n2333, Z => 
                           n4982);
   U2611 : AO4 port map( A => n4010, B => n1367, C => n2443, D => n2332, Z => 
                           n4983);
   U2612 : AO4 port map( A => n4011, B => n1411, C => n2443, D => n2331, Z => 
                           n4984);
   U2613 : AO4 port map( A => n4008, B => n575, C => n362, D => n2330, Z => 
                           n4985);
   U2614 : AO4 port map( A => n4009, B => n619, C => n2443, D => n2329, Z => 
                           n4986);
   U2615 : AO4 port map( A => n4006, B => n663, C => n2443, D => n2328, Z => 
                           n4987);
   U2616 : AO4 port map( A => n4007, B => n707, C => n362, D => n2327, Z => 
                           n4988);
   U2617 : AO4 port map( A => n4092, B => n390, C => n361, D => n2382, Z => 
                           n5509);
   U2618 : AO4 port map( A => n4093, B => n399, C => n2452, D => n2381, Z => 
                           n5510);
   U2619 : AO4 port map( A => n4090, B => n400, C => n361, D => n2380, Z => 
                           n5511);
   U2620 : AO4 port map( A => n4091, B => n401, C => n2452, D => n2379, Z => 
                           n5512);
   U2621 : AO4 port map( A => n4088, B => n402, C => n361, D => n2378, Z => 
                           n5513);
   U2622 : AO4 port map( A => n4089, B => n403, C => n2452, D => n2377, Z => 
                           n5514);
   U2623 : AO4 port map( A => n4086, B => n404, C => n361, D => n2376, Z => 
                           n5515);
   U2624 : AO4 port map( A => n4087, B => n405, C => n2452, D => n2375, Z => 
                           n5516);
   U2625 : AO4 port map( A => n4100, B => n406, C => n361, D => n2374, Z => 
                           n5517);
   U2626 : AO4 port map( A => n4101, B => n411, C => n2452, D => n2373, Z => 
                           n5518);
   U2627 : AO4 port map( A => n4098, B => n412, C => n2452, D => n2372, Z => 
                           n5519);
   U2628 : AO4 port map( A => n4099, B => n413, C => n2452, D => n2371, Z => 
                           n5520);
   U2629 : AO4 port map( A => n4096, B => n414, C => n2452, D => n2370, Z => 
                           n5521);
   U2630 : AO4 port map( A => n4097, B => n415, C => n2452, D => n2369, Z => 
                           n5522);
   U2631 : AO4 port map( A => n4094, B => n416, C => n361, D => n2368, Z => 
                           n5523);
   U2632 : AO4 port map( A => n4095, B => n417, C => n2452, D => n2367, Z => 
                           n5524);
   U2633 : AO4 port map( A => n4108, B => n418, C => n2452, D => n2366, Z => 
                           n5525);
   U2634 : AO4 port map( A => n4109, B => n423, C => n361, D => n2365, Z => 
                           n5526);
   U2635 : AO4 port map( A => n4106, B => n424, C => n2452, D => n2364, Z => 
                           n5527);
   U2636 : AO4 port map( A => n4107, B => n425, C => n2452, D => n2363, Z => 
                           n5528);
   U2637 : AO4 port map( A => n4104, B => n426, C => n361, D => n2362, Z => 
                           n5529);
   U2638 : AO4 port map( A => n4105, B => n427, C => n2452, D => n2361, Z => 
                           n5530);
   U2639 : AO4 port map( A => n4102, B => n428, C => n2452, D => n2360, Z => 
                           n5531);
   U2640 : AO4 port map( A => n4103, B => n429, C => n361, D => n2359, Z => 
                           n5532);
   U2641 : AO4 port map( A => n4052, B => n751, C => n2452, D => n2358, Z => 
                           n5533);
   U2642 : AO4 port map( A => n4053, B => n795, C => n2452, D => n2357, Z => 
                           n5534);
   U2643 : AO4 port map( A => n4050, B => n839, C => n361, D => n2356, Z => 
                           n5535);
   U2644 : AO4 port map( A => n4051, B => n883, C => n2452, D => n2355, Z => 
                           n5536);
   U2645 : AO4 port map( A => n4048, B => n430, C => n361, D => n2354, Z => 
                           n5537);
   U2646 : AO4 port map( A => n4049, B => n435, C => n361, D => n2353, Z => 
                           n5538);
   U2647 : AO4 port map( A => n4046, B => n436, C => n361, D => n2352, Z => 
                           n5539);
   U2648 : AO4 port map( A => n4047, B => n437, C => n361, D => n2351, Z => 
                           n5540);
   U2649 : AO4 port map( A => n4060, B => n927, C => n361, D => n2350, Z => 
                           n5541);
   U2650 : AO4 port map( A => n4061, B => n971, C => n361, D => n2349, Z => 
                           n5542);
   U2651 : AO4 port map( A => n4058, B => n1015, C => n361, D => n2348, Z => 
                           n5543);
   U2652 : AO4 port map( A => n4059, B => n1059, C => n361, D => n2347, Z => 
                           n5544);
   U2653 : AO4 port map( A => n4056, B => n438, C => n361, D => n2346, Z => 
                           n5545);
   U2654 : AO4 port map( A => n4057, B => n439, C => n361, D => n2345, Z => 
                           n5546);
   U2655 : AO4 port map( A => n4054, B => n440, C => n361, D => n2344, Z => 
                           n5547);
   U2656 : AO4 port map( A => n4055, B => n441, C => n361, D => n2343, Z => 
                           n5548);
   U2657 : AO4 port map( A => n4068, B => n1103, C => n361, D => n2342, Z => 
                           n5549);
   U2658 : AO4 port map( A => n4069, B => n1147, C => n361, D => n2341, Z => 
                           n5550);
   U2659 : AO4 port map( A => n4066, B => n1191, C => n361, D => n2340, Z => 
                           n5551);
   U2660 : AO4 port map( A => n4067, B => n1235, C => n361, D => n2339, Z => 
                           n5552);
   U2661 : AO4 port map( A => n4064, B => n442, C => n361, D => n2338, Z => 
                           n5553);
   U2662 : AO4 port map( A => n4065, B => n443, C => n361, D => n2337, Z => 
                           n5554);
   U2663 : AO4 port map( A => n4062, B => n487, C => n361, D => n2336, Z => 
                           n5555);
   U2664 : AO4 port map( A => n4063, B => n531, C => n2452, D => n2335, Z => 
                           n5556);
   U2665 : AO4 port map( A => n4076, B => n1279, C => n2452, D => n2334, Z => 
                           n5557);
   U2666 : AO4 port map( A => n4077, B => n1323, C => n2452, D => n2333, Z => 
                           n5558);
   U2667 : AO4 port map( A => n4074, B => n1367, C => n2452, D => n2332, Z => 
                           n5559);
   U2668 : AO4 port map( A => n4075, B => n1411, C => n2452, D => n2331, Z => 
                           n5560);
   U2669 : AO4 port map( A => n4072, B => n575, C => n2452, D => n2330, Z => 
                           n5561);
   U2670 : AO4 port map( A => n4073, B => n619, C => n2452, D => n2329, Z => 
                           n5562);
   U2671 : AO4 port map( A => n4070, B => n663, C => n2452, D => n2328, Z => 
                           n5563);
   U2672 : AO4 port map( A => n4071, B => n707, C => n2452, D => n2327, Z => 
                           n5564);
   U2673 : AO4 port map( A => n4156, B => n390, C => n293, D => n2382, Z => 
                           n6021);
   U2674 : AO4 port map( A => n4157, B => n399, C => n293, D => n2381, Z => 
                           n6022);
   U2675 : AO4 port map( A => n4154, B => n400, C => n293, D => n2380, Z => 
                           n6023);
   U2676 : AO4 port map( A => n4155, B => n401, C => n2460, D => n2379, Z => 
                           n6024);
   U2677 : AO4 port map( A => n4152, B => n402, C => n2460, D => n2378, Z => 
                           n6025);
   U2678 : AO4 port map( A => n4153, B => n403, C => n2460, D => n2377, Z => 
                           n6026);
   U2679 : AO4 port map( A => n4150, B => n404, C => n2460, D => n2376, Z => 
                           n6027);
   U2680 : AO4 port map( A => n4151, B => n405, C => n2460, D => n2375, Z => 
                           n6028);
   U2681 : AO4 port map( A => n4164, B => n406, C => n2460, D => n2374, Z => 
                           n6029);
   U2682 : AO4 port map( A => n4165, B => n411, C => n2460, D => n2373, Z => 
                           n6030);
   U2683 : AO4 port map( A => n4162, B => n412, C => n2460, D => n2372, Z => 
                           n6031);
   U2684 : AO4 port map( A => n4163, B => n413, C => n2460, D => n2371, Z => 
                           n6032);
   U2685 : AO4 port map( A => n4160, B => n414, C => n2460, D => n2370, Z => 
                           n6033);
   U2686 : AO4 port map( A => n4161, B => n415, C => n2460, D => n2369, Z => 
                           n6034);
   U2687 : AO4 port map( A => n4158, B => n416, C => n293, D => n2368, Z => 
                           n6035);
   U2688 : AO4 port map( A => n4159, B => n417, C => n2460, D => n2367, Z => 
                           n6036);
   U2689 : AO4 port map( A => n4172, B => n418, C => n293, D => n2366, Z => 
                           n6037);
   U2690 : AO4 port map( A => n4173, B => n423, C => n2460, D => n2365, Z => 
                           n6038);
   U2691 : AO4 port map( A => n4170, B => n424, C => n293, D => n2364, Z => 
                           n6039);
   U2692 : AO4 port map( A => n4171, B => n425, C => n2460, D => n2363, Z => 
                           n6040);
   U2693 : AO4 port map( A => n4168, B => n426, C => n293, D => n2362, Z => 
                           n6041);
   U2694 : AO4 port map( A => n4169, B => n427, C => n2460, D => n2361, Z => 
                           n6042);
   U2695 : AO4 port map( A => n4166, B => n428, C => n2460, D => n2360, Z => 
                           n6043);
   U2696 : AO4 port map( A => n4167, B => n429, C => n2460, D => n2359, Z => 
                           n6044);
   U2697 : AO4 port map( A => n4116, B => n751, C => n2460, D => n2358, Z => 
                           n6045);
   U2698 : AO4 port map( A => n4117, B => n795, C => n2460, D => n2357, Z => 
                           n6046);
   U2699 : AO4 port map( A => n4114, B => n839, C => n2460, D => n2356, Z => 
                           n6047);
   U2700 : AO4 port map( A => n4115, B => n883, C => n2460, D => n2355, Z => 
                           n6048);
   U2701 : AO4 port map( A => n4112, B => n430, C => n293, D => n2354, Z => 
                           n6049);
   U2702 : AO4 port map( A => n4113, B => n435, C => n2460, D => n2353, Z => 
                           n6050);
   U2703 : AO4 port map( A => n4110, B => n436, C => n2460, D => n2352, Z => 
                           n6051);
   U2704 : AO4 port map( A => n4111, B => n437, C => n293, D => n2351, Z => 
                           n6052);
   U2705 : AO4 port map( A => n4124, B => n927, C => n2460, D => n2350, Z => 
                           n6053);
   U2706 : AO4 port map( A => n4125, B => n971, C => n2460, D => n2349, Z => 
                           n6054);
   U2707 : AO4 port map( A => n4122, B => n1015, C => n293, D => n2348, Z => 
                           n6055);
   U2708 : AO4 port map( A => n4123, B => n1059, C => n293, D => n2347, Z => 
                           n6056);
   U2709 : AO4 port map( A => n4120, B => n438, C => n293, D => n2346, Z => 
                           n6057);
   U2710 : AO4 port map( A => n4121, B => n439, C => n293, D => n2345, Z => 
                           n6058);
   U2711 : AO4 port map( A => n4118, B => n440, C => n293, D => n2344, Z => 
                           n6059);
   U2712 : AO4 port map( A => n4119, B => n441, C => n293, D => n2343, Z => 
                           n6060);
   U2713 : AO4 port map( A => n4132, B => n1103, C => n2460, D => n2342, Z => 
                           n6061);
   U2714 : AO4 port map( A => n4133, B => n1147, C => n2460, D => n2341, Z => 
                           n6062);
   U2715 : AO4 port map( A => n4130, B => n1191, C => n293, D => n2340, Z => 
                           n6063);
   U2716 : AO4 port map( A => n4131, B => n1235, C => n293, D => n2339, Z => 
                           n6064);
   U2717 : AO4 port map( A => n4128, B => n442, C => n293, D => n2338, Z => 
                           n6065);
   U2718 : AO4 port map( A => n4129, B => n443, C => n293, D => n2337, Z => 
                           n6066);
   U2719 : AO4 port map( A => n4126, B => n487, C => n293, D => n2336, Z => 
                           n6067);
   U2720 : AO4 port map( A => n4127, B => n531, C => n293, D => n2335, Z => 
                           n6068);
   U2721 : AO4 port map( A => n4140, B => n1279, C => n293, D => n2334, Z => 
                           n6069);
   U2722 : AO4 port map( A => n4141, B => n1323, C => n293, D => n2333, Z => 
                           n6070);
   U2723 : AO4 port map( A => n4138, B => n1367, C => n293, D => n2332, Z => 
                           n6071);
   U2724 : AO4 port map( A => n4139, B => n1411, C => n293, D => n2331, Z => 
                           n6072);
   U2725 : AO4 port map( A => n4136, B => n575, C => n293, D => n2330, Z => 
                           n6073);
   U2726 : AO4 port map( A => n4137, B => n619, C => n293, D => n2329, Z => 
                           n6074);
   U2727 : AO4 port map( A => n4134, B => n663, C => n293, D => n2328, Z => 
                           n6075);
   U2728 : AO4 port map( A => n4135, B => n707, C => n293, D => n2327, Z => 
                           n6076);
   U2729 : AO4 port map( A => n4220, B => n390, C => n286, D => n2382, Z => 
                           n6533);
   U2730 : AO4 port map( A => n4221, B => n399, C => n2468, D => n2381, Z => 
                           n6534);
   U2731 : AO4 port map( A => n4218, B => n400, C => n286, D => n2380, Z => 
                           n6535);
   U2732 : AO4 port map( A => n4219, B => n401, C => n2468, D => n2379, Z => 
                           n6536);
   U2733 : AO4 port map( A => n4216, B => n402, C => n286, D => n2378, Z => 
                           n6537);
   U2734 : AO4 port map( A => n4217, B => n403, C => n2468, D => n2377, Z => 
                           n6538);
   U2735 : AO4 port map( A => n4214, B => n404, C => n286, D => n2376, Z => 
                           n6539);
   U2736 : AO4 port map( A => n4215, B => n405, C => n2468, D => n2375, Z => 
                           n6540);
   U2737 : AO4 port map( A => n4228, B => n406, C => n286, D => n2374, Z => 
                           n6541);
   U2738 : AO4 port map( A => n4229, B => n411, C => n2468, D => n2373, Z => 
                           n6542);
   U2739 : AO4 port map( A => n4226, B => n412, C => n2468, D => n2372, Z => 
                           n6543);
   U2740 : AO4 port map( A => n4227, B => n413, C => n2468, D => n2371, Z => 
                           n6544);
   U2741 : AO4 port map( A => n4224, B => n414, C => n2468, D => n2370, Z => 
                           n6545);
   U2742 : AO4 port map( A => n4225, B => n415, C => n2468, D => n2369, Z => 
                           n6546);
   U2743 : AO4 port map( A => n4222, B => n416, C => n286, D => n2368, Z => 
                           n6547);
   U2744 : AO4 port map( A => n4223, B => n417, C => n2468, D => n2367, Z => 
                           n6548);
   U2745 : AO4 port map( A => n4236, B => n418, C => n2468, D => n2366, Z => 
                           n6549);
   U2746 : AO4 port map( A => n4237, B => n423, C => n286, D => n2365, Z => 
                           n6550);
   U2747 : AO4 port map( A => n4234, B => n424, C => n2468, D => n2364, Z => 
                           n6551);
   U2748 : AO4 port map( A => n4235, B => n425, C => n2468, D => n2363, Z => 
                           n6552);
   U2749 : AO4 port map( A => n4232, B => n426, C => n286, D => n2362, Z => 
                           n6553);
   U2750 : AO4 port map( A => n4233, B => n427, C => n2468, D => n2361, Z => 
                           n6554);
   U2751 : AO4 port map( A => n4230, B => n428, C => n2468, D => n2360, Z => 
                           n6555);
   U2752 : AO4 port map( A => n4231, B => n429, C => n286, D => n2359, Z => 
                           n6556);
   U2753 : AO4 port map( A => n4180, B => n751, C => n2468, D => n2358, Z => 
                           n6557);
   U2754 : AO4 port map( A => n4181, B => n795, C => n2468, D => n2357, Z => 
                           n6558);
   U2755 : AO4 port map( A => n4178, B => n839, C => n286, D => n2356, Z => 
                           n6559);
   U2756 : AO4 port map( A => n4179, B => n883, C => n2468, D => n2355, Z => 
                           n6560);
   U2757 : AO4 port map( A => n4176, B => n430, C => n286, D => n2354, Z => 
                           n6561);
   U2758 : AO4 port map( A => n4177, B => n435, C => n286, D => n2353, Z => 
                           n6562);
   U2759 : AO4 port map( A => n4174, B => n436, C => n286, D => n2352, Z => 
                           n6563);
   U2760 : AO4 port map( A => n4175, B => n437, C => n286, D => n2351, Z => 
                           n6564);
   U2761 : AO4 port map( A => n4188, B => n927, C => n286, D => n2350, Z => 
                           n6565);
   U2762 : AO4 port map( A => n4189, B => n971, C => n286, D => n2349, Z => 
                           n6566);
   U2763 : AO4 port map( A => n4186, B => n1015, C => n286, D => n2348, Z => 
                           n6567);
   U2764 : AO4 port map( A => n4187, B => n1059, C => n286, D => n2347, Z => 
                           n6568);
   U2765 : AO4 port map( A => n4184, B => n438, C => n286, D => n2346, Z => 
                           n6569);
   U2766 : AO4 port map( A => n4185, B => n439, C => n286, D => n2345, Z => 
                           n6570);
   U2767 : AO4 port map( A => n4182, B => n440, C => n286, D => n2344, Z => 
                           n6571);
   U2768 : AO4 port map( A => n4183, B => n441, C => n286, D => n2343, Z => 
                           n6572);
   U2769 : AO4 port map( A => n4196, B => n1103, C => n286, D => n2342, Z => 
                           n6573);
   U2770 : AO4 port map( A => n4197, B => n1147, C => n286, D => n2341, Z => 
                           n6574);
   U2771 : AO4 port map( A => n4194, B => n1191, C => n286, D => n2340, Z => 
                           n6575);
   U2772 : AO4 port map( A => n4195, B => n1235, C => n286, D => n2339, Z => 
                           n6576);
   U2773 : AO4 port map( A => n4192, B => n442, C => n286, D => n2338, Z => 
                           n6577);
   U2774 : AO4 port map( A => n4193, B => n443, C => n286, D => n2337, Z => 
                           n6578);
   U2775 : AO4 port map( A => n4190, B => n487, C => n286, D => n2336, Z => 
                           n6579);
   U2776 : AO4 port map( A => n4191, B => n531, C => n2468, D => n2335, Z => 
                           n6580);
   U2777 : AO4 port map( A => n4204, B => n1279, C => n2468, D => n2334, Z => 
                           n6581);
   U2778 : AO4 port map( A => n4205, B => n1323, C => n2468, D => n2333, Z => 
                           n6582);
   U2779 : AO4 port map( A => n4202, B => n1367, C => n2468, D => n2332, Z => 
                           n6583);
   U2780 : AO4 port map( A => n4203, B => n1411, C => n2468, D => n2331, Z => 
                           n6584);
   U2781 : AO4 port map( A => n4200, B => n575, C => n2468, D => n2330, Z => 
                           n6585);
   U2782 : AO4 port map( A => n4201, B => n619, C => n2468, D => n2329, Z => 
                           n6586);
   U2783 : AO4 port map( A => n4198, B => n663, C => n2468, D => n2328, Z => 
                           n6587);
   U2784 : AO4 port map( A => n4199, B => n707, C => n2468, D => n2327, Z => 
                           n6588);
   U2785 : AO4 port map( A => n4284, B => n390, C => n360, D => n2382, Z => 
                           n4997);
   U2786 : AO4 port map( A => n4285, B => n399, C => n360, D => n2381, Z => 
                           n4998);
   U2787 : AO4 port map( A => n4282, B => n400, C => n360, D => n2380, Z => 
                           n4999);
   U2788 : AO4 port map( A => n4283, B => n401, C => n2444, D => n2379, Z => 
                           n5000);
   U2789 : AO4 port map( A => n4280, B => n402, C => n2444, D => n2378, Z => 
                           n5001);
   U2790 : AO4 port map( A => n4281, B => n403, C => n2444, D => n2377, Z => 
                           n5002);
   U2791 : AO4 port map( A => n4278, B => n404, C => n2444, D => n2376, Z => 
                           n5003);
   U2792 : AO4 port map( A => n4279, B => n405, C => n2444, D => n2375, Z => 
                           n5004);
   U2793 : AO4 port map( A => n4292, B => n406, C => n2444, D => n2374, Z => 
                           n5005);
   U2794 : AO4 port map( A => n4293, B => n411, C => n2444, D => n2373, Z => 
                           n5006);
   U2795 : AO4 port map( A => n4290, B => n412, C => n2444, D => n2372, Z => 
                           n5007);
   U2796 : AO4 port map( A => n4291, B => n413, C => n2444, D => n2371, Z => 
                           n5008);
   U2797 : AO4 port map( A => n4288, B => n414, C => n2444, D => n2370, Z => 
                           n5009);
   U2798 : AO4 port map( A => n4289, B => n415, C => n2444, D => n2369, Z => 
                           n5010);
   U2799 : AO4 port map( A => n4286, B => n416, C => n360, D => n2368, Z => 
                           n5011);
   U2800 : AO4 port map( A => n4287, B => n417, C => n2444, D => n2367, Z => 
                           n5012);
   U2801 : AO4 port map( A => n4300, B => n418, C => n360, D => n2366, Z => 
                           n5013);
   U2802 : AO4 port map( A => n4301, B => n423, C => n2444, D => n2365, Z => 
                           n5014);
   U2803 : AO4 port map( A => n4298, B => n424, C => n360, D => n2364, Z => 
                           n5015);
   U2804 : AO4 port map( A => n4299, B => n425, C => n2444, D => n2363, Z => 
                           n5016);
   U2805 : AO4 port map( A => n4296, B => n426, C => n360, D => n2362, Z => 
                           n5017);
   U2806 : AO4 port map( A => n4297, B => n427, C => n2444, D => n2361, Z => 
                           n5018);
   U2807 : AO4 port map( A => n4294, B => n428, C => n2444, D => n2360, Z => 
                           n5019);
   U2808 : AO4 port map( A => n4295, B => n429, C => n2444, D => n2359, Z => 
                           n5020);
   U2809 : AO4 port map( A => n4244, B => n751, C => n2444, D => n2358, Z => 
                           n5021);
   U2810 : AO4 port map( A => n4245, B => n795, C => n2444, D => n2357, Z => 
                           n5022);
   U2811 : AO4 port map( A => n4242, B => n839, C => n2444, D => n2356, Z => 
                           n5023);
   U2812 : AO4 port map( A => n4243, B => n883, C => n2444, D => n2355, Z => 
                           n5024);
   U2813 : AO4 port map( A => n4240, B => n430, C => n360, D => n2354, Z => 
                           n5025);
   U2814 : AO4 port map( A => n4241, B => n435, C => n2444, D => n2353, Z => 
                           n5026);
   U2815 : AO4 port map( A => n4238, B => n436, C => n2444, D => n2352, Z => 
                           n5027);
   U2816 : AO4 port map( A => n4239, B => n437, C => n360, D => n2351, Z => 
                           n5028);
   U2817 : AO4 port map( A => n4252, B => n927, C => n2444, D => n2350, Z => 
                           n5029);
   U2818 : AO4 port map( A => n4253, B => n971, C => n2444, D => n2349, Z => 
                           n5030);
   U2819 : AO4 port map( A => n4250, B => n1015, C => n360, D => n2348, Z => 
                           n5031);
   U2820 : AO4 port map( A => n4251, B => n1059, C => n360, D => n2347, Z => 
                           n5032);
   U2821 : AO4 port map( A => n4248, B => n438, C => n360, D => n2346, Z => 
                           n5033);
   U2822 : AO4 port map( A => n4249, B => n439, C => n360, D => n2345, Z => 
                           n5034);
   U2823 : AO4 port map( A => n4246, B => n440, C => n360, D => n2344, Z => 
                           n5035);
   U2824 : AO4 port map( A => n4247, B => n441, C => n360, D => n2343, Z => 
                           n5036);
   U2825 : AO4 port map( A => n4260, B => n1103, C => n2444, D => n2342, Z => 
                           n5037);
   U2826 : AO4 port map( A => n4261, B => n1147, C => n2444, D => n2341, Z => 
                           n5038);
   U2827 : AO4 port map( A => n4258, B => n1191, C => n360, D => n2340, Z => 
                           n5039);
   U2828 : AO4 port map( A => n4259, B => n1235, C => n360, D => n2339, Z => 
                           n5040);
   U2829 : AO4 port map( A => n4256, B => n442, C => n360, D => n2338, Z => 
                           n5041);
   U2830 : AO4 port map( A => n4257, B => n443, C => n360, D => n2337, Z => 
                           n5042);
   U2831 : AO4 port map( A => n4254, B => n487, C => n360, D => n2336, Z => 
                           n5043);
   U2832 : AO4 port map( A => n4255, B => n531, C => n360, D => n2335, Z => 
                           n5044);
   U2833 : AO4 port map( A => n4268, B => n1279, C => n360, D => n2334, Z => 
                           n5045);
   U2834 : AO4 port map( A => n4269, B => n1323, C => n360, D => n2333, Z => 
                           n5046);
   U2835 : AO4 port map( A => n4266, B => n1367, C => n360, D => n2332, Z => 
                           n5047);
   U2836 : AO4 port map( A => n4267, B => n1411, C => n360, D => n2331, Z => 
                           n5048);
   U2837 : AO4 port map( A => n4264, B => n575, C => n360, D => n2330, Z => 
                           n5049);
   U2838 : AO4 port map( A => n4265, B => n619, C => n360, D => n2329, Z => 
                           n5050);
   U2839 : AO4 port map( A => n4262, B => n663, C => n360, D => n2328, Z => 
                           n5051);
   U2840 : AO4 port map( A => n4263, B => n707, C => n360, D => n2327, Z => 
                           n5052);
   U2841 : AO4 port map( A => n4348, B => n390, C => n359, D => n2382, Z => 
                           n5573);
   U2842 : AO4 port map( A => n4349, B => n399, C => n2453, D => n2381, Z => 
                           n5574);
   U2843 : AO4 port map( A => n4346, B => n400, C => n359, D => n2380, Z => 
                           n5575);
   U2844 : AO4 port map( A => n4347, B => n401, C => n2453, D => n2379, Z => 
                           n5576);
   U2845 : AO4 port map( A => n4344, B => n402, C => n359, D => n2378, Z => 
                           n5577);
   U2846 : AO4 port map( A => n4345, B => n403, C => n2453, D => n2377, Z => 
                           n5578);
   U2847 : AO4 port map( A => n4342, B => n404, C => n359, D => n2376, Z => 
                           n5579);
   U2848 : AO4 port map( A => n4343, B => n405, C => n2453, D => n2375, Z => 
                           n5580);
   U2849 : AO4 port map( A => n4356, B => n406, C => n359, D => n2374, Z => 
                           n5581);
   U2850 : AO4 port map( A => n4357, B => n411, C => n2453, D => n2373, Z => 
                           n5582);
   U2851 : AO4 port map( A => n4354, B => n412, C => n2453, D => n2372, Z => 
                           n5583);
   U2852 : AO4 port map( A => n4355, B => n413, C => n2453, D => n2371, Z => 
                           n5584);
   U2853 : AO4 port map( A => n4352, B => n414, C => n2453, D => n2370, Z => 
                           n5585);
   U2854 : AO4 port map( A => n4353, B => n415, C => n2453, D => n2369, Z => 
                           n5586);
   U2855 : AO4 port map( A => n4350, B => n416, C => n359, D => n2368, Z => 
                           n5587);
   U2856 : AO4 port map( A => n4351, B => n417, C => n2453, D => n2367, Z => 
                           n5588);
   U2857 : AO4 port map( A => n4364, B => n418, C => n2453, D => n2366, Z => 
                           n5589);
   U2858 : AO4 port map( A => n4365, B => n423, C => n359, D => n2365, Z => 
                           n5590);
   U2859 : AO4 port map( A => n4362, B => n424, C => n2453, D => n2364, Z => 
                           n5591);
   U2860 : AO4 port map( A => n4363, B => n425, C => n2453, D => n2363, Z => 
                           n5592);
   U2861 : AO4 port map( A => n4360, B => n426, C => n359, D => n2362, Z => 
                           n5593);
   U2862 : AO4 port map( A => n4361, B => n427, C => n2453, D => n2361, Z => 
                           n5594);
   U2863 : AO4 port map( A => n4358, B => n428, C => n2453, D => n2360, Z => 
                           n5595);
   U2864 : AO4 port map( A => n4359, B => n429, C => n359, D => n2359, Z => 
                           n5596);
   U2865 : AO4 port map( A => n4308, B => n751, C => n2453, D => n2358, Z => 
                           n5597);
   U2866 : AO4 port map( A => n4309, B => n795, C => n2453, D => n2357, Z => 
                           n5598);
   U2867 : AO4 port map( A => n4306, B => n839, C => n359, D => n2356, Z => 
                           n5599);
   U2868 : AO4 port map( A => n4307, B => n883, C => n2453, D => n2355, Z => 
                           n5600);
   U2869 : AO4 port map( A => n4304, B => n430, C => n359, D => n2354, Z => 
                           n5601);
   U2870 : AO4 port map( A => n4305, B => n435, C => n359, D => n2353, Z => 
                           n5602);
   U2871 : AO4 port map( A => n4302, B => n436, C => n359, D => n2352, Z => 
                           n5603);
   U2872 : AO4 port map( A => n4303, B => n437, C => n359, D => n2351, Z => 
                           n5604);
   U2873 : AO4 port map( A => n4316, B => n927, C => n359, D => n2350, Z => 
                           n5605);
   U2874 : AO4 port map( A => n4317, B => n971, C => n359, D => n2349, Z => 
                           n5606);
   U2875 : AO4 port map( A => n4314, B => n1015, C => n359, D => n2348, Z => 
                           n5607);
   U2876 : AO4 port map( A => n4315, B => n1059, C => n359, D => n2347, Z => 
                           n5608);
   U2877 : AO4 port map( A => n4312, B => n438, C => n359, D => n2346, Z => 
                           n5609);
   U2878 : AO4 port map( A => n4313, B => n439, C => n359, D => n2345, Z => 
                           n5610);
   U2879 : AO4 port map( A => n4310, B => n440, C => n359, D => n2344, Z => 
                           n5611);
   U2880 : AO4 port map( A => n4311, B => n441, C => n359, D => n2343, Z => 
                           n5612);
   U2881 : AO4 port map( A => n4324, B => n1103, C => n359, D => n2342, Z => 
                           n5613);
   U2882 : AO4 port map( A => n4325, B => n1147, C => n359, D => n2341, Z => 
                           n5614);
   U2883 : AO4 port map( A => n4322, B => n1191, C => n359, D => n2340, Z => 
                           n5615);
   U2884 : AO4 port map( A => n4323, B => n1235, C => n359, D => n2339, Z => 
                           n5616);
   U2885 : AO4 port map( A => n4320, B => n442, C => n359, D => n2338, Z => 
                           n5617);
   U2886 : AO4 port map( A => n4321, B => n443, C => n359, D => n2337, Z => 
                           n5618);
   U2887 : AO4 port map( A => n4318, B => n487, C => n359, D => n2336, Z => 
                           n5619);
   U2888 : AO4 port map( A => n4319, B => n531, C => n2453, D => n2335, Z => 
                           n5620);
   U2889 : AO4 port map( A => n4332, B => n1279, C => n2453, D => n2334, Z => 
                           n5621);
   U2890 : AO4 port map( A => n4333, B => n1323, C => n2453, D => n2333, Z => 
                           n5622);
   U2891 : AO4 port map( A => n4330, B => n1367, C => n2453, D => n2332, Z => 
                           n5623);
   U2892 : AO4 port map( A => n4331, B => n1411, C => n2453, D => n2331, Z => 
                           n5624);
   U2893 : AO4 port map( A => n4328, B => n575, C => n2453, D => n2330, Z => 
                           n5625);
   U2894 : AO4 port map( A => n4329, B => n619, C => n2453, D => n2329, Z => 
                           n5626);
   U2895 : AO4 port map( A => n4326, B => n663, C => n2453, D => n2328, Z => 
                           n5627);
   U2896 : AO4 port map( A => n4327, B => n707, C => n2453, D => n2327, Z => 
                           n5628);
   U2897 : AO4 port map( A => n4412, B => n390, C => n284, D => n2382, Z => 
                           n6085);
   U2898 : AO4 port map( A => n4413, B => n399, C => n2461, D => n2381, Z => 
                           n6086);
   U2899 : AO4 port map( A => n4410, B => n400, C => n284, D => n2380, Z => 
                           n6087);
   U2900 : AO4 port map( A => n4411, B => n401, C => n2461, D => n2379, Z => 
                           n6088);
   U2901 : AO4 port map( A => n4408, B => n402, C => n284, D => n2378, Z => 
                           n6089);
   U2902 : AO4 port map( A => n4409, B => n403, C => n2461, D => n2377, Z => 
                           n6090);
   U2903 : AO4 port map( A => n4406, B => n404, C => n284, D => n2376, Z => 
                           n6091);
   U2904 : AO4 port map( A => n4407, B => n405, C => n2461, D => n2375, Z => 
                           n6092);
   U2905 : AO4 port map( A => n4420, B => n406, C => n284, D => n2374, Z => 
                           n6093);
   U2906 : AO4 port map( A => n4421, B => n411, C => n2461, D => n2373, Z => 
                           n6094);
   U2907 : AO4 port map( A => n4418, B => n412, C => n2461, D => n2372, Z => 
                           n6095);
   U2908 : AO4 port map( A => n4419, B => n413, C => n2461, D => n2371, Z => 
                           n6096);
   U2909 : AO4 port map( A => n4416, B => n414, C => n2461, D => n2370, Z => 
                           n6097);
   U2910 : AO4 port map( A => n4417, B => n415, C => n2461, D => n2369, Z => 
                           n6098);
   U2911 : AO4 port map( A => n4414, B => n416, C => n284, D => n2368, Z => 
                           n6099);
   U2912 : AO4 port map( A => n4415, B => n417, C => n2461, D => n2367, Z => 
                           n6100);
   U2913 : AO4 port map( A => n4428, B => n418, C => n2461, D => n2366, Z => 
                           n6101);
   U2914 : AO4 port map( A => n4429, B => n423, C => n284, D => n2365, Z => 
                           n6102);
   U2915 : AO4 port map( A => n4426, B => n424, C => n2461, D => n2364, Z => 
                           n6103);
   U2916 : AO4 port map( A => n4427, B => n425, C => n2461, D => n2363, Z => 
                           n6104);
   U2917 : AO4 port map( A => n4424, B => n426, C => n284, D => n2362, Z => 
                           n6105);
   U2918 : AO4 port map( A => n4425, B => n427, C => n2461, D => n2361, Z => 
                           n6106);
   U2919 : AO4 port map( A => n4422, B => n428, C => n2461, D => n2360, Z => 
                           n6107);
   U2920 : AO4 port map( A => n4423, B => n429, C => n284, D => n2359, Z => 
                           n6108);
   U2921 : AO4 port map( A => n4372, B => n751, C => n2461, D => n2358, Z => 
                           n6109);
   U2922 : AO4 port map( A => n4373, B => n795, C => n2461, D => n2357, Z => 
                           n6110);
   U2923 : AO4 port map( A => n4370, B => n839, C => n284, D => n2356, Z => 
                           n6111);
   U2924 : AO4 port map( A => n4371, B => n883, C => n2461, D => n2355, Z => 
                           n6112);
   U2925 : AO4 port map( A => n4368, B => n430, C => n284, D => n2354, Z => 
                           n6113);
   U2926 : AO4 port map( A => n4369, B => n435, C => n284, D => n2353, Z => 
                           n6114);
   U2927 : AO4 port map( A => n4366, B => n436, C => n284, D => n2352, Z => 
                           n6115);
   U2928 : AO4 port map( A => n4367, B => n437, C => n284, D => n2351, Z => 
                           n6116);
   U2929 : AO4 port map( A => n4380, B => n927, C => n284, D => n2350, Z => 
                           n6117);
   U2930 : AO4 port map( A => n4381, B => n971, C => n284, D => n2349, Z => 
                           n6118);
   U2931 : AO4 port map( A => n4378, B => n1015, C => n284, D => n2348, Z => 
                           n6119);
   U2932 : AO4 port map( A => n4379, B => n1059, C => n284, D => n2347, Z => 
                           n6120);
   U2933 : AO4 port map( A => n4376, B => n438, C => n284, D => n2346, Z => 
                           n6121);
   U2934 : AO4 port map( A => n4377, B => n439, C => n284, D => n2345, Z => 
                           n6122);
   U2935 : AO4 port map( A => n4374, B => n440, C => n284, D => n2344, Z => 
                           n6123);
   U2936 : AO4 port map( A => n4375, B => n441, C => n284, D => n2343, Z => 
                           n6124);
   U2937 : AO4 port map( A => n4388, B => n1103, C => n284, D => n2342, Z => 
                           n6125);
   U2938 : AO4 port map( A => n4389, B => n1147, C => n284, D => n2341, Z => 
                           n6126);
   U2939 : AO4 port map( A => n4386, B => n1191, C => n284, D => n2340, Z => 
                           n6127);
   U2940 : AO4 port map( A => n4387, B => n1235, C => n284, D => n2339, Z => 
                           n6128);
   U2941 : AO4 port map( A => n4384, B => n442, C => n284, D => n2338, Z => 
                           n6129);
   U2942 : AO4 port map( A => n4385, B => n443, C => n284, D => n2337, Z => 
                           n6130);
   U2943 : AO4 port map( A => n4382, B => n487, C => n284, D => n2336, Z => 
                           n6131);
   U2944 : AO4 port map( A => n4383, B => n531, C => n2461, D => n2335, Z => 
                           n6132);
   U2945 : AO4 port map( A => n4396, B => n1279, C => n2461, D => n2334, Z => 
                           n6133);
   U2946 : AO4 port map( A => n4397, B => n1323, C => n2461, D => n2333, Z => 
                           n6134);
   U2947 : AO4 port map( A => n4394, B => n1367, C => n2461, D => n2332, Z => 
                           n6135);
   U2948 : AO4 port map( A => n4395, B => n1411, C => n2461, D => n2331, Z => 
                           n6136);
   U2949 : AO4 port map( A => n4392, B => n575, C => n2461, D => n2330, Z => 
                           n6137);
   U2950 : AO4 port map( A => n4393, B => n619, C => n2461, D => n2329, Z => 
                           n6138);
   U2951 : AO4 port map( A => n4390, B => n663, C => n2461, D => n2328, Z => 
                           n6139);
   U2952 : AO4 port map( A => n4391, B => n707, C => n2461, D => n2327, Z => 
                           n6140);
   U2953 : AO4 port map( A => n4476, B => n390, C => n2469, D => n2382, Z => 
                           n6597);
   U2954 : AO4 port map( A => n4477, B => n399, C => n2469, D => n2381, Z => 
                           n6598);
   U2955 : AO4 port map( A => n4474, B => n400, C => n2469, D => n2380, Z => 
                           n6599);
   U2956 : AO4 port map( A => n4475, B => n401, C => n2469, D => n2379, Z => 
                           n6600);
   U2957 : AO4 port map( A => n4472, B => n402, C => n2469, D => n2378, Z => 
                           n6601);
   U2958 : AO4 port map( A => n4473, B => n403, C => n2469, D => n2377, Z => 
                           n6602);
   U2959 : AO4 port map( A => n4470, B => n404, C => n2469, D => n2376, Z => 
                           n6603);
   U2960 : AO4 port map( A => n4471, B => n405, C => n2469, D => n2375, Z => 
                           n6604);
   U2961 : AO4 port map( A => n4484, B => n406, C => n276, D => n2374, Z => 
                           n6605);
   U2962 : AO4 port map( A => n4485, B => n411, C => n2469, D => n2373, Z => 
                           n6606);
   U2963 : AO4 port map( A => n4482, B => n412, C => n2469, D => n2372, Z => 
                           n6607);
   U2964 : AO4 port map( A => n4483, B => n413, C => n2469, D => n2371, Z => 
                           n6608);
   U2965 : AO4 port map( A => n4480, B => n414, C => n276, D => n2370, Z => 
                           n6609);
   U2966 : AO4 port map( A => n4481, B => n415, C => n2469, D => n2369, Z => 
                           n6610);
   U2967 : AO4 port map( A => n4478, B => n416, C => n276, D => n2368, Z => 
                           n6611);
   U2968 : AO4 port map( A => n4479, B => n417, C => n276, D => n2367, Z => 
                           n6612);
   U2969 : AO4 port map( A => n4492, B => n418, C => n276, D => n2366, Z => 
                           n6613);
   U2970 : AO4 port map( A => n4493, B => n423, C => n276, D => n2365, Z => 
                           n6614);
   U2971 : AO4 port map( A => n4490, B => n424, C => n276, D => n2364, Z => 
                           n6615);
   U2972 : AO4 port map( A => n4491, B => n425, C => n276, D => n2363, Z => 
                           n6616);
   U2973 : AO4 port map( A => n4488, B => n426, C => n276, D => n2362, Z => 
                           n6617);
   U2974 : AO4 port map( A => n4489, B => n427, C => n276, D => n2361, Z => 
                           n6618);
   U2975 : AO4 port map( A => n4486, B => n428, C => n276, D => n2360, Z => 
                           n6619);
   U2976 : AO4 port map( A => n4487, B => n429, C => n276, D => n2359, Z => 
                           n6620);
   U2977 : AO4 port map( A => n4436, B => n751, C => n276, D => n2358, Z => 
                           n6621);
   U2978 : AO4 port map( A => n4437, B => n795, C => n276, D => n2357, Z => 
                           n6622);
   U2979 : AO4 port map( A => n4434, B => n839, C => n276, D => n2356, Z => 
                           n6623);
   U2980 : AO4 port map( A => n4435, B => n883, C => n276, D => n2355, Z => 
                           n6624);
   U2981 : AO4 port map( A => n4432, B => n430, C => n276, D => n2354, Z => 
                           n6625);
   U2982 : AO4 port map( A => n4433, B => n435, C => n276, D => n2353, Z => 
                           n6626);
   U2983 : AO4 port map( A => n4430, B => n436, C => n276, D => n2352, Z => 
                           n6627);
   U2984 : AO4 port map( A => n4431, B => n437, C => n276, D => n2351, Z => 
                           n6628);
   U2985 : AO4 port map( A => n4444, B => n927, C => n276, D => n2350, Z => 
                           n6629);
   U2986 : AO4 port map( A => n4445, B => n971, C => n276, D => n2349, Z => 
                           n6630);
   U2987 : AO4 port map( A => n4442, B => n1015, C => n276, D => n2348, Z => 
                           n6631);
   U2988 : AO4 port map( A => n4443, B => n1059, C => n276, D => n2347, Z => 
                           n6632);
   U2989 : AO4 port map( A => n4440, B => n438, C => n276, D => n2346, Z => 
                           n6633);
   U2990 : AO4 port map( A => n4441, B => n439, C => n276, D => n2345, Z => 
                           n6634);
   U2991 : AO4 port map( A => n4438, B => n440, C => n2469, D => n2344, Z => 
                           n6635);
   U2992 : AO4 port map( A => n4439, B => n441, C => n2469, D => n2343, Z => 
                           n6636);
   U2993 : AO4 port map( A => n4452, B => n1103, C => n2469, D => n2342, Z => 
                           n6637);
   U2994 : AO4 port map( A => n4453, B => n1147, C => n2469, D => n2341, Z => 
                           n6638);
   U2995 : AO4 port map( A => n4450, B => n1191, C => n2469, D => n2340, Z => 
                           n6639);
   U2996 : AO4 port map( A => n4451, B => n1235, C => n276, D => n2339, Z => 
                           n6640);
   U2997 : AO4 port map( A => n4448, B => n442, C => n2469, D => n2338, Z => 
                           n6641);
   U2998 : AO4 port map( A => n4449, B => n443, C => n2469, D => n2337, Z => 
                           n6642);
   U2999 : AO4 port map( A => n4446, B => n487, C => n276, D => n2336, Z => 
                           n6643);
   U3000 : AO4 port map( A => n4447, B => n531, C => n2469, D => n2335, Z => 
                           n6644);
   U3001 : AO4 port map( A => n4460, B => n1279, C => n2469, D => n2334, Z => 
                           n6645);
   U3002 : AO4 port map( A => n4461, B => n1323, C => n276, D => n2333, Z => 
                           n6646);
   U3003 : AO4 port map( A => n4458, B => n1367, C => n2469, D => n2332, Z => 
                           n6647);
   U3004 : AO4 port map( A => n4459, B => n1411, C => n2469, D => n2331, Z => 
                           n6648);
   U3005 : AO4 port map( A => n4456, B => n575, C => n276, D => n2330, Z => 
                           n6649);
   U3006 : AO4 port map( A => n4457, B => n619, C => n2469, D => n2329, Z => 
                           n6650);
   U3007 : AO4 port map( A => n4454, B => n663, C => n2469, D => n2328, Z => 
                           n6651);
   U3008 : AO4 port map( A => n4455, B => n707, C => n276, D => n2327, Z => 
                           n6652);
   U3009 : AO4 port map( A => n4540, B => n390, C => n354, D => n2382, Z => 
                           n5061);
   U3010 : AO4 port map( A => n4541, B => n399, C => n2445, D => n2381, Z => 
                           n5062);
   U3011 : AO4 port map( A => n4538, B => n400, C => n354, D => n2380, Z => 
                           n5063);
   U3012 : AO4 port map( A => n4539, B => n401, C => n2445, D => n2379, Z => 
                           n5064);
   U3013 : AO4 port map( A => n4536, B => n402, C => n354, D => n2378, Z => 
                           n5065);
   U3014 : AO4 port map( A => n4537, B => n403, C => n2445, D => n2377, Z => 
                           n5066);
   U3015 : AO4 port map( A => n4534, B => n404, C => n354, D => n2376, Z => 
                           n5067);
   U3016 : AO4 port map( A => n4535, B => n405, C => n2445, D => n2375, Z => 
                           n5068);
   U3017 : AO4 port map( A => n4548, B => n406, C => n354, D => n2374, Z => 
                           n5069);
   U3018 : AO4 port map( A => n4549, B => n411, C => n2445, D => n2373, Z => 
                           n5070);
   U3019 : AO4 port map( A => n4546, B => n412, C => n2445, D => n2372, Z => 
                           n5071);
   U3020 : AO4 port map( A => n4547, B => n413, C => n2445, D => n2371, Z => 
                           n5072);
   U3021 : AO4 port map( A => n4544, B => n414, C => n2445, D => n2370, Z => 
                           n5073);
   U3022 : AO4 port map( A => n4545, B => n415, C => n2445, D => n2369, Z => 
                           n5074);
   U3023 : AO4 port map( A => n4542, B => n416, C => n354, D => n2368, Z => 
                           n5075);
   U3024 : AO4 port map( A => n4543, B => n417, C => n2445, D => n2367, Z => 
                           n5076);
   U3025 : AO4 port map( A => n4556, B => n418, C => n2445, D => n2366, Z => 
                           n5077);
   U3026 : AO4 port map( A => n4557, B => n423, C => n354, D => n2365, Z => 
                           n5078);
   U3027 : AO4 port map( A => n4554, B => n424, C => n2445, D => n2364, Z => 
                           n5079);
   U3028 : AO4 port map( A => n4555, B => n425, C => n2445, D => n2363, Z => 
                           n5080);
   U3029 : AO4 port map( A => n4552, B => n426, C => n354, D => n2362, Z => 
                           n5081);
   U3030 : AO4 port map( A => n4553, B => n427, C => n2445, D => n2361, Z => 
                           n5082);
   U3031 : AO4 port map( A => n4550, B => n428, C => n2445, D => n2360, Z => 
                           n5083);
   U3032 : AO4 port map( A => n4551, B => n429, C => n354, D => n2359, Z => 
                           n5084);
   U3033 : AO4 port map( A => n4500, B => n751, C => n2445, D => n2358, Z => 
                           n5085);
   U3034 : AO4 port map( A => n4501, B => n795, C => n2445, D => n2357, Z => 
                           n5086);
   U3035 : AO4 port map( A => n4498, B => n839, C => n354, D => n2356, Z => 
                           n5087);
   U3036 : AO4 port map( A => n4499, B => n883, C => n2445, D => n2355, Z => 
                           n5088);
   U3037 : AO4 port map( A => n4496, B => n430, C => n354, D => n2354, Z => 
                           n5089);
   U3038 : AO4 port map( A => n4497, B => n435, C => n354, D => n2353, Z => 
                           n5090);
   U3039 : AO4 port map( A => n4494, B => n436, C => n354, D => n2352, Z => 
                           n5091);
   U3040 : AO4 port map( A => n4495, B => n437, C => n354, D => n2351, Z => 
                           n5092);
   U3041 : AO4 port map( A => n4508, B => n927, C => n354, D => n2350, Z => 
                           n5093);
   U3042 : AO4 port map( A => n4509, B => n971, C => n354, D => n2349, Z => 
                           n5094);
   U3043 : AO4 port map( A => n4506, B => n1015, C => n354, D => n2348, Z => 
                           n5095);
   U3044 : AO4 port map( A => n4507, B => n1059, C => n354, D => n2347, Z => 
                           n5096);
   U3045 : AO4 port map( A => n4504, B => n438, C => n354, D => n2346, Z => 
                           n5097);
   U3046 : AO4 port map( A => n4505, B => n439, C => n354, D => n2345, Z => 
                           n5098);
   U3047 : AO4 port map( A => n4502, B => n440, C => n354, D => n2344, Z => 
                           n5099);
   U3048 : AO4 port map( A => n4503, B => n441, C => n354, D => n2343, Z => 
                           n5100);
   U3049 : AO4 port map( A => n4516, B => n1103, C => n354, D => n2342, Z => 
                           n5101);
   U3050 : AO4 port map( A => n4517, B => n1147, C => n354, D => n2341, Z => 
                           n5102);
   U3051 : AO4 port map( A => n4514, B => n1191, C => n354, D => n2340, Z => 
                           n5103);
   U3052 : AO4 port map( A => n4515, B => n1235, C => n354, D => n2339, Z => 
                           n5104);
   U3053 : AO4 port map( A => n4512, B => n442, C => n354, D => n2338, Z => 
                           n5105);
   U3054 : AO4 port map( A => n4513, B => n443, C => n354, D => n2337, Z => 
                           n5106);
   U3055 : AO4 port map( A => n4510, B => n487, C => n354, D => n2336, Z => 
                           n5107);
   U3056 : AO4 port map( A => n4511, B => n531, C => n2445, D => n2335, Z => 
                           n5108);
   U3057 : AO4 port map( A => n4524, B => n1279, C => n2445, D => n2334, Z => 
                           n5109);
   U3058 : AO4 port map( A => n4525, B => n1323, C => n2445, D => n2333, Z => 
                           n5110);
   U3059 : AO4 port map( A => n4522, B => n1367, C => n2445, D => n2332, Z => 
                           n5111);
   U3060 : AO4 port map( A => n4523, B => n1411, C => n2445, D => n2331, Z => 
                           n5112);
   U3061 : AO4 port map( A => n4520, B => n575, C => n2445, D => n2330, Z => 
                           n5113);
   U3062 : AO4 port map( A => n4521, B => n619, C => n2445, D => n2329, Z => 
                           n5114);
   U3063 : AO4 port map( A => n4518, B => n663, C => n2445, D => n2328, Z => 
                           n5115);
   U3064 : AO4 port map( A => n4519, B => n707, C => n2445, D => n2327, Z => 
                           n5116);
   U3065 : NR4 port map( A => n343, B => n344, C => n345, D => n346, Z => n342)
                           ;
   U3066 : AO4 port map( A => n2543, B => n81, C => n2542, D => n229, Z => n343
                           );
   U3067 : AO4 port map( A => n2545, B => n270, C => n2544, D => n272, Z => 
                           n344);
   U3068 : AO4 port map( A => n2547, B => n72, C => n2546, D => n228, Z => n345
                           );
   U3069 : NR4 port map( A => n355, B => n356, C => n357, D => n358, Z => n341)
                           ;
   U3070 : AO4 port map( A => n2551, B => n71, C => n2550, D => n227, Z => n355
                           );
   U3071 : AO4 port map( A => n2553, B => n255, C => n2552, D => n257, Z => 
                           n356);
   U3072 : AO4 port map( A => n2555, B => n12, C => n2554, D => n23, Z => n357)
                           ;
   U3073 : NR4 port map( A => n367, B => n368, C => n369, D => n370, Z => n340)
                           ;
   U3074 : AO4 port map( A => n2559, B => n69, C => n2558, D => n224, Z => n367
                           );
   U3075 : AO4 port map( A => n2561, B => n265, C => n2560, D => n269, Z => 
                           n368);
   U3076 : AO4 port map( A => n2563, B => n11, C => n2562, D => n217, Z => n369
                           );
   U3077 : NR4 port map( A => n379, B => n380, C => n381, D => n382, Z => n339)
                           ;
   U3078 : AO4 port map( A => n2567, B => n59, C => n2566, D => n209, Z => n379
                           );
   U3079 : AO4 port map( A => n2569, B => n251, C => n2568, D => n253, Z => 
                           n380);
   U3080 : AO4 port map( A => n2571, B => n10, C => n2570, D => n22, Z => n381)
                           ;
   U3081 : NR4 port map( A => n395, B => n396, C => n397, D => n398, Z => n394)
                           ;
   U3082 : AO4 port map( A => n2511, B => n58, C => n2510, D => n200, Z => n395
                           );
   U3083 : AO4 port map( A => n2513, B => n260, C => n2512, D => n261, Z => 
                           n396);
   U3084 : AO4 port map( A => n2515, B => n9, C => n2514, D => n180, Z => n397)
                           ;
   U3085 : NR4 port map( A => n407, B => n408, C => n409, D => n410, Z => n393)
                           ;
   U3086 : AO4 port map( A => n2519, B => n53, C => n2518, D => n170, Z => n407
                           );
   U3087 : AO4 port map( A => n2521, B => n249, C => n2520, D => n250, Z => 
                           n408);
   U3088 : AO4 port map( A => n2523, B => n28, C => n2522, D => n14, Z => n409)
                           ;
   U3089 : NR4 port map( A => n419, B => n420, C => n421, D => n422, Z => n392)
                           ;
   U3090 : AO4 port map( A => n2527, B => n8, C => n2526, D => n163, Z => n419)
                           ;
   U3091 : AO4 port map( A => n2529, B => n258, C => n2528, D => n259, Z => 
                           n420);
   U3092 : AO4 port map( A => n2531, B => n7, C => n2530, D => n150, Z => n421)
                           ;
   U3093 : NR4 port map( A => n431, B => n432, C => n433, D => n434, Z => n391)
                           ;
   U3094 : AO4 port map( A => n2535, B => n48, C => n2534, D => n122, Z => n431
                           );
   U3095 : AO4 port map( A => n2537, B => n246, C => n2536, D => n248, Z => 
                           n432);
   U3096 : AO4 port map( A => n2539, B => n6, C => n2538, D => n109, Z => n433)
                           ;
   U3097 : NR4 port map( A => n451, B => n452, C => n453, D => n454, Z => n450)
                           ;
   U3098 : AO4 port map( A => n2607, B => n81, C => n2606, D => n229, Z => n451
                           );
   U3099 : AO4 port map( A => n2609, B => n270, C => n2608, D => n272, Z => 
                           n452);
   U3100 : AO4 port map( A => n2611, B => n72, C => n2610, D => n228, Z => n453
                           );
   U3101 : NR4 port map( A => n455, B => n456, C => n457, D => n458, Z => n449)
                           ;
   U3102 : AO4 port map( A => n2615, B => n71, C => n2614, D => n227, Z => n455
                           );
   U3103 : AO4 port map( A => n2617, B => n255, C => n2616, D => n257, Z => 
                           n456);
   U3104 : AO4 port map( A => n2619, B => n12, C => n2618, D => n23, Z => n457)
                           ;
   U3105 : NR4 port map( A => n459, B => n460, C => n461, D => n462, Z => n448)
                           ;
   U3106 : AO4 port map( A => n2623, B => n69, C => n2622, D => n224, Z => n459
                           );
   U3107 : AO4 port map( A => n2625, B => n265, C => n2624, D => n269, Z => 
                           n460);
   U3108 : AO4 port map( A => n2627, B => n11, C => n2626, D => n217, Z => n461
                           );
   U3109 : NR4 port map( A => n463, B => n464, C => n465, D => n466, Z => n447)
                           ;
   U3110 : AO4 port map( A => n2631, B => n59, C => n2630, D => n209, Z => n463
                           );
   U3111 : AO4 port map( A => n2633, B => n251, C => n2632, D => n253, Z => 
                           n464);
   U3112 : AO4 port map( A => n2635, B => n10, C => n2634, D => n22, Z => n465)
                           ;
   U3113 : NR4 port map( A => n471, B => n472, C => n473, D => n474, Z => n470)
                           ;
   U3114 : AO4 port map( A => n2575, B => n58, C => n2574, D => n200, Z => n471
                           );
   U3115 : AO4 port map( A => n2577, B => n260, C => n2576, D => n261, Z => 
                           n472);
   U3116 : AO4 port map( A => n2579, B => n9, C => n2578, D => n180, Z => n473)
                           ;
   U3117 : NR4 port map( A => n475, B => n476, C => n477, D => n478, Z => n469)
                           ;
   U3118 : AO4 port map( A => n2583, B => n53, C => n2582, D => n170, Z => n475
                           );
   U3119 : AO4 port map( A => n2585, B => n249, C => n2584, D => n250, Z => 
                           n476);
   U3120 : AO4 port map( A => n2587, B => n28, C => n2586, D => n14, Z => n477)
                           ;
   U3121 : NR4 port map( A => n479, B => n480, C => n481, D => n482, Z => n468)
                           ;
   U3122 : AO4 port map( A => n2591, B => n8, C => n2590, D => n163, Z => n479)
                           ;
   U3123 : AO4 port map( A => n2593, B => n258, C => n2592, D => n259, Z => 
                           n480);
   U3124 : AO4 port map( A => n2595, B => n7, C => n2594, D => n150, Z => n481)
                           ;
   U3125 : NR4 port map( A => n483, B => n484, C => n485, D => n486, Z => n467)
                           ;
   U3126 : AO4 port map( A => n2599, B => n48, C => n2598, D => n122, Z => n483
                           );
   U3127 : AO4 port map( A => n2601, B => n246, C => n2600, D => n248, Z => 
                           n484);
   U3128 : AO4 port map( A => n2603, B => n6, C => n2602, D => n109, Z => n485)
                           ;
   U3129 : NR4 port map( A => n495, B => n496, C => n497, D => n498, Z => n494)
                           ;
   U3130 : AO4 port map( A => n2671, B => n81, C => n2670, D => n229, Z => n495
                           );
   U3131 : AO4 port map( A => n2673, B => n270, C => n2672, D => n272, Z => 
                           n496);
   U3132 : AO4 port map( A => n2675, B => n72, C => n2674, D => n228, Z => n497
                           );
   U3133 : NR4 port map( A => n499, B => n500, C => n501, D => n502, Z => n493)
                           ;
   U3134 : AO4 port map( A => n2679, B => n71, C => n2678, D => n227, Z => n499
                           );
   U3135 : AO4 port map( A => n2681, B => n255, C => n2680, D => n257, Z => 
                           n500);
   U3136 : AO4 port map( A => n2683, B => n12, C => n2682, D => n23, Z => n501)
                           ;
   U3137 : NR4 port map( A => n503, B => n504, C => n505, D => n506, Z => n492)
                           ;
   U3138 : AO4 port map( A => n2687, B => n69, C => n2686, D => n224, Z => n503
                           );
   U3139 : AO4 port map( A => n2689, B => n265, C => n2688, D => n269, Z => 
                           n504);
   U3140 : AO4 port map( A => n2691, B => n11, C => n2690, D => n217, Z => n505
                           );
   U3141 : NR4 port map( A => n507, B => n508, C => n509, D => n510, Z => n491)
                           ;
   U3142 : AO4 port map( A => n2695, B => n59, C => n2694, D => n209, Z => n507
                           );
   U3143 : AO4 port map( A => n2697, B => n251, C => n2696, D => n253, Z => 
                           n508);
   U3144 : AO4 port map( A => n2699, B => n10, C => n2698, D => n22, Z => n509)
                           ;
   U3145 : NR4 port map( A => n515, B => n516, C => n517, D => n518, Z => n514)
                           ;
   U3146 : AO4 port map( A => n2639, B => n58, C => n2638, D => n200, Z => n515
                           );
   U3147 : AO4 port map( A => n2641, B => n260, C => n2640, D => n261, Z => 
                           n516);
   U3148 : AO4 port map( A => n2643, B => n9, C => n2642, D => n180, Z => n517)
                           ;
   U3149 : NR4 port map( A => n519, B => n520, C => n521, D => n522, Z => n513)
                           ;
   U3150 : AO4 port map( A => n2647, B => n53, C => n2646, D => n170, Z => n519
                           );
   U3151 : AO4 port map( A => n2649, B => n249, C => n2648, D => n250, Z => 
                           n520);
   U3152 : AO4 port map( A => n2651, B => n28, C => n2650, D => n14, Z => n521)
                           ;
   U3153 : NR4 port map( A => n523, B => n524, C => n525, D => n526, Z => n512)
                           ;
   U3154 : AO4 port map( A => n2655, B => n8, C => n2654, D => n163, Z => n523)
                           ;
   U3155 : AO4 port map( A => n2657, B => n258, C => n2656, D => n259, Z => 
                           n524);
   U3156 : AO4 port map( A => n2659, B => n7, C => n2658, D => n150, Z => n525)
                           ;
   U3157 : NR4 port map( A => n527, B => n528, C => n529, D => n530, Z => n511)
                           ;
   U3158 : AO4 port map( A => n2663, B => n48, C => n2662, D => n122, Z => n527
                           );
   U3159 : AO4 port map( A => n2665, B => n246, C => n2664, D => n248, Z => 
                           n528);
   U3160 : AO4 port map( A => n2667, B => n6, C => n2666, D => n109, Z => n529)
                           ;
   U3161 : NR4 port map( A => n539, B => n540, C => n541, D => n542, Z => n538)
                           ;
   U3162 : AO4 port map( A => n2735, B => n81, C => n2734, D => n229, Z => n539
                           );
   U3163 : AO4 port map( A => n2737, B => n270, C => n2736, D => n272, Z => 
                           n540);
   U3164 : AO4 port map( A => n2739, B => n72, C => n2738, D => n228, Z => n541
                           );
   U3165 : NR4 port map( A => n543, B => n544, C => n545, D => n546, Z => n537)
                           ;
   U3166 : AO4 port map( A => n2743, B => n71, C => n2742, D => n227, Z => n543
                           );
   U3167 : AO4 port map( A => n2745, B => n255, C => n2744, D => n257, Z => 
                           n544);
   U3168 : AO4 port map( A => n2747, B => n12, C => n2746, D => n23, Z => n545)
                           ;
   U3169 : NR4 port map( A => n547, B => n548, C => n549, D => n550, Z => n536)
                           ;
   U3170 : AO4 port map( A => n2751, B => n69, C => n2750, D => n224, Z => n547
                           );
   U3171 : AO4 port map( A => n2753, B => n265, C => n2752, D => n269, Z => 
                           n548);
   U3172 : AO4 port map( A => n2755, B => n11, C => n2754, D => n217, Z => n549
                           );
   U3173 : NR4 port map( A => n551, B => n552, C => n553, D => n554, Z => n535)
                           ;
   U3174 : AO4 port map( A => n2759, B => n59, C => n2758, D => n209, Z => n551
                           );
   U3175 : AO4 port map( A => n2761, B => n251, C => n2760, D => n253, Z => 
                           n552);
   U3176 : AO4 port map( A => n2763, B => n10, C => n2762, D => n22, Z => n553)
                           ;
   U3177 : NR4 port map( A => n559, B => n560, C => n561, D => n562, Z => n558)
                           ;
   U3178 : AO4 port map( A => n2703, B => n58, C => n2702, D => n200, Z => n559
                           );
   U3179 : AO4 port map( A => n2705, B => n260, C => n2704, D => n261, Z => 
                           n560);
   U3180 : AO4 port map( A => n2707, B => n9, C => n2706, D => n180, Z => n561)
                           ;
   U3181 : NR4 port map( A => n563, B => n564, C => n565, D => n566, Z => n557)
                           ;
   U3182 : AO4 port map( A => n2711, B => n53, C => n2710, D => n170, Z => n563
                           );
   U3183 : AO4 port map( A => n2713, B => n249, C => n2712, D => n250, Z => 
                           n564);
   U3184 : AO4 port map( A => n2715, B => n28, C => n2714, D => n14, Z => n565)
                           ;
   U3185 : NR4 port map( A => n567, B => n568, C => n569, D => n570, Z => n556)
                           ;
   U3186 : AO4 port map( A => n2719, B => n8, C => n2718, D => n163, Z => n567)
                           ;
   U3187 : AO4 port map( A => n2721, B => n258, C => n2720, D => n259, Z => 
                           n568);
   U3188 : AO4 port map( A => n2723, B => n7, C => n2722, D => n150, Z => n569)
                           ;
   U3189 : NR4 port map( A => n571, B => n572, C => n573, D => n574, Z => n555)
                           ;
   U3190 : AO4 port map( A => n2727, B => n48, C => n2726, D => n122, Z => n571
                           );
   U3191 : AO4 port map( A => n2729, B => n246, C => n2728, D => n248, Z => 
                           n572);
   U3192 : AO4 port map( A => n2731, B => n6, C => n2730, D => n109, Z => n573)
                           ;
   U3193 : NR4 port map( A => n583, B => n584, C => n585, D => n586, Z => n582)
                           ;
   U3194 : AO4 port map( A => n2799, B => n81, C => n2798, D => n229, Z => n583
                           );
   U3195 : AO4 port map( A => n2801, B => n270, C => n2800, D => n272, Z => 
                           n584);
   U3196 : AO4 port map( A => n2803, B => n72, C => n2802, D => n228, Z => n585
                           );
   U3197 : NR4 port map( A => n587, B => n588, C => n589, D => n590, Z => n581)
                           ;
   U3198 : AO4 port map( A => n2807, B => n71, C => n2806, D => n227, Z => n587
                           );
   U3199 : AO4 port map( A => n2809, B => n255, C => n2808, D => n257, Z => 
                           n588);
   U3200 : AO4 port map( A => n2811, B => n12, C => n2810, D => n23, Z => n589)
                           ;
   U3201 : NR4 port map( A => n591, B => n592, C => n593, D => n594, Z => n580)
                           ;
   U3202 : AO4 port map( A => n2815, B => n69, C => n2814, D => n224, Z => n591
                           );
   U3203 : AO4 port map( A => n2817, B => n265, C => n2816, D => n269, Z => 
                           n592);
   U3204 : AO4 port map( A => n2819, B => n11, C => n2818, D => n217, Z => n593
                           );
   U3205 : NR4 port map( A => n595, B => n596, C => n597, D => n598, Z => n579)
                           ;
   U3206 : AO4 port map( A => n2823, B => n59, C => n2822, D => n209, Z => n595
                           );
   U3207 : AO4 port map( A => n2825, B => n251, C => n2824, D => n253, Z => 
                           n596);
   U3208 : AO4 port map( A => n2827, B => n10, C => n2826, D => n22, Z => n597)
                           ;
   U3209 : NR4 port map( A => n603, B => n604, C => n605, D => n606, Z => n602)
                           ;
   U3210 : AO4 port map( A => n2767, B => n58, C => n2766, D => n200, Z => n603
                           );
   U3211 : AO4 port map( A => n2769, B => n260, C => n2768, D => n261, Z => 
                           n604);
   U3212 : AO4 port map( A => n2771, B => n9, C => n2770, D => n180, Z => n605)
                           ;
   U3213 : NR4 port map( A => n607, B => n608, C => n609, D => n610, Z => n601)
                           ;
   U3214 : AO4 port map( A => n2775, B => n53, C => n2774, D => n170, Z => n607
                           );
   U3215 : AO4 port map( A => n2777, B => n249, C => n2776, D => n250, Z => 
                           n608);
   U3216 : AO4 port map( A => n2779, B => n28, C => n2778, D => n14, Z => n609)
                           ;
   U3217 : NR4 port map( A => n611, B => n612, C => n613, D => n614, Z => n600)
                           ;
   U3218 : AO4 port map( A => n2783, B => n8, C => n2782, D => n163, Z => n611)
                           ;
   U3219 : AO4 port map( A => n2785, B => n258, C => n2784, D => n259, Z => 
                           n612);
   U3220 : AO4 port map( A => n2787, B => n7, C => n2786, D => n150, Z => n613)
                           ;
   U3221 : NR4 port map( A => n615, B => n616, C => n617, D => n618, Z => n599)
                           ;
   U3222 : AO4 port map( A => n2791, B => n48, C => n2790, D => n122, Z => n615
                           );
   U3223 : AO4 port map( A => n2793, B => n246, C => n2792, D => n248, Z => 
                           n616);
   U3224 : AO4 port map( A => n2795, B => n6, C => n2794, D => n109, Z => n617)
                           ;
   U3225 : NR4 port map( A => n627, B => n628, C => n629, D => n630, Z => n626)
                           ;
   U3226 : AO4 port map( A => n2863, B => n81, C => n2862, D => n229, Z => n627
                           );
   U3227 : AO4 port map( A => n2865, B => n270, C => n2864, D => n272, Z => 
                           n628);
   U3228 : AO4 port map( A => n2867, B => n72, C => n2866, D => n228, Z => n629
                           );
   U3229 : NR4 port map( A => n631, B => n632, C => n633, D => n634, Z => n625)
                           ;
   U3230 : AO4 port map( A => n2871, B => n71, C => n2870, D => n227, Z => n631
                           );
   U3231 : AO4 port map( A => n2873, B => n255, C => n2872, D => n257, Z => 
                           n632);
   U3232 : AO4 port map( A => n2875, B => n12, C => n2874, D => n23, Z => n633)
                           ;
   U3233 : NR4 port map( A => n635, B => n636, C => n637, D => n638, Z => n624)
                           ;
   U3234 : AO4 port map( A => n2879, B => n69, C => n2878, D => n224, Z => n635
                           );
   U3235 : AO4 port map( A => n2881, B => n265, C => n2880, D => n269, Z => 
                           n636);
   U3236 : AO4 port map( A => n2883, B => n11, C => n2882, D => n217, Z => n637
                           );
   U3237 : NR4 port map( A => n639, B => n640, C => n641, D => n642, Z => n623)
                           ;
   U3238 : AO4 port map( A => n2887, B => n59, C => n2886, D => n209, Z => n639
                           );
   U3239 : AO4 port map( A => n2889, B => n251, C => n2888, D => n253, Z => 
                           n640);
   U3240 : AO4 port map( A => n2891, B => n10, C => n2890, D => n22, Z => n641)
                           ;
   U3241 : NR4 port map( A => n647, B => n648, C => n649, D => n650, Z => n646)
                           ;
   U3242 : AO4 port map( A => n2831, B => n58, C => n2830, D => n200, Z => n647
                           );
   U3243 : AO4 port map( A => n2833, B => n260, C => n2832, D => n261, Z => 
                           n648);
   U3244 : AO4 port map( A => n2835, B => n9, C => n2834, D => n180, Z => n649)
                           ;
   U3245 : NR4 port map( A => n651, B => n652, C => n653, D => n654, Z => n645)
                           ;
   U3246 : AO4 port map( A => n2839, B => n53, C => n2838, D => n170, Z => n651
                           );
   U3247 : AO4 port map( A => n2841, B => n249, C => n2840, D => n250, Z => 
                           n652);
   U3248 : AO4 port map( A => n2843, B => n28, C => n2842, D => n14, Z => n653)
                           ;
   U3249 : NR4 port map( A => n655, B => n656, C => n657, D => n658, Z => n644)
                           ;
   U3250 : AO4 port map( A => n2847, B => n8, C => n2846, D => n163, Z => n655)
                           ;
   U3251 : AO4 port map( A => n2849, B => n258, C => n2848, D => n259, Z => 
                           n656);
   U3252 : AO4 port map( A => n2851, B => n7, C => n2850, D => n150, Z => n657)
                           ;
   U3253 : NR4 port map( A => n659, B => n660, C => n661, D => n662, Z => n643)
                           ;
   U3254 : AO4 port map( A => n2855, B => n48, C => n2854, D => n122, Z => n659
                           );
   U3255 : AO4 port map( A => n2857, B => n246, C => n2856, D => n248, Z => 
                           n660);
   U3256 : AO4 port map( A => n2859, B => n6, C => n2858, D => n109, Z => n661)
                           ;
   U3257 : NR4 port map( A => n671, B => n672, C => n673, D => n674, Z => n670)
                           ;
   U3258 : AO4 port map( A => n2927, B => n81, C => n2926, D => n229, Z => n671
                           );
   U3259 : AO4 port map( A => n2929, B => n270, C => n2928, D => n272, Z => 
                           n672);
   U3260 : AO4 port map( A => n2931, B => n72, C => n2930, D => n228, Z => n673
                           );
   U3261 : NR4 port map( A => n675, B => n676, C => n677, D => n678, Z => n669)
                           ;
   U3262 : AO4 port map( A => n2935, B => n71, C => n2934, D => n227, Z => n675
                           );
   U3263 : AO4 port map( A => n2937, B => n255, C => n2936, D => n257, Z => 
                           n676);
   U3264 : AO4 port map( A => n2939, B => n12, C => n2938, D => n23, Z => n677)
                           ;
   U3265 : NR4 port map( A => n679, B => n680, C => n681, D => n682, Z => n668)
                           ;
   U3266 : AO4 port map( A => n2943, B => n69, C => n2942, D => n224, Z => n679
                           );
   U3267 : AO4 port map( A => n2945, B => n265, C => n2944, D => n269, Z => 
                           n680);
   U3268 : AO4 port map( A => n2947, B => n11, C => n2946, D => n217, Z => n681
                           );
   U3269 : NR4 port map( A => n683, B => n684, C => n685, D => n686, Z => n667)
                           ;
   U3270 : AO4 port map( A => n2951, B => n59, C => n2950, D => n209, Z => n683
                           );
   U3271 : AO4 port map( A => n2953, B => n251, C => n2952, D => n253, Z => 
                           n684);
   U3272 : AO4 port map( A => n2955, B => n10, C => n2954, D => n22, Z => n685)
                           ;
   U3273 : NR4 port map( A => n691, B => n692, C => n693, D => n694, Z => n690)
                           ;
   U3274 : AO4 port map( A => n2895, B => n58, C => n2894, D => n200, Z => n691
                           );
   U3275 : AO4 port map( A => n2897, B => n260, C => n2896, D => n261, Z => 
                           n692);
   U3276 : AO4 port map( A => n2899, B => n9, C => n2898, D => n180, Z => n693)
                           ;
   U3277 : NR4 port map( A => n695, B => n696, C => n697, D => n698, Z => n689)
                           ;
   U3278 : AO4 port map( A => n2903, B => n53, C => n2902, D => n170, Z => n695
                           );
   U3279 : AO4 port map( A => n2905, B => n249, C => n2904, D => n250, Z => 
                           n696);
   U3280 : AO4 port map( A => n2907, B => n28, C => n2906, D => n14, Z => n697)
                           ;
   U3281 : NR4 port map( A => n699, B => n700, C => n701, D => n702, Z => n688)
                           ;
   U3282 : AO4 port map( A => n2911, B => n8, C => n2910, D => n163, Z => n699)
                           ;
   U3283 : AO4 port map( A => n2913, B => n258, C => n2912, D => n259, Z => 
                           n700);
   U3284 : AO4 port map( A => n2915, B => n7, C => n2914, D => n150, Z => n701)
                           ;
   U3285 : NR4 port map( A => n703, B => n704, C => n705, D => n706, Z => n687)
                           ;
   U3286 : AO4 port map( A => n2919, B => n48, C => n2918, D => n122, Z => n703
                           );
   U3287 : AO4 port map( A => n2921, B => n246, C => n2920, D => n248, Z => 
                           n704);
   U3288 : AO4 port map( A => n2923, B => n6, C => n2922, D => n109, Z => n705)
                           ;
   U3289 : NR4 port map( A => n715, B => n716, C => n717, D => n718, Z => n714)
                           ;
   U3290 : AO4 port map( A => n2991, B => n81, C => n2990, D => n229, Z => n715
                           );
   U3291 : AO4 port map( A => n2993, B => n270, C => n2992, D => n272, Z => 
                           n716);
   U3292 : AO4 port map( A => n2995, B => n72, C => n2994, D => n228, Z => n717
                           );
   U3293 : NR4 port map( A => n719, B => n720, C => n721, D => n722, Z => n713)
                           ;
   U3294 : AO4 port map( A => n2999, B => n71, C => n2998, D => n227, Z => n719
                           );
   U3295 : AO4 port map( A => n3001, B => n255, C => n3000, D => n257, Z => 
                           n720);
   U3296 : AO4 port map( A => n3003, B => n12, C => n3002, D => n23, Z => n721)
                           ;
   U3297 : NR4 port map( A => n723, B => n724, C => n725, D => n726, Z => n712)
                           ;
   U3298 : AO4 port map( A => n3007, B => n69, C => n3006, D => n224, Z => n723
                           );
   U3299 : AO4 port map( A => n3009, B => n265, C => n3008, D => n269, Z => 
                           n724);
   U3300 : AO4 port map( A => n3011, B => n11, C => n3010, D => n217, Z => n725
                           );
   U3301 : NR4 port map( A => n727, B => n728, C => n729, D => n730, Z => n711)
                           ;
   U3302 : AO4 port map( A => n3015, B => n59, C => n3014, D => n209, Z => n727
                           );
   U3303 : AO4 port map( A => n3017, B => n251, C => n3016, D => n253, Z => 
                           n728);
   U3304 : AO4 port map( A => n3019, B => n10, C => n3018, D => n22, Z => n729)
                           ;
   U3305 : NR4 port map( A => n735, B => n736, C => n737, D => n738, Z => n734)
                           ;
   U3306 : AO4 port map( A => n2959, B => n58, C => n2958, D => n200, Z => n735
                           );
   U3307 : AO4 port map( A => n2961, B => n260, C => n2960, D => n261, Z => 
                           n736);
   U3308 : AO4 port map( A => n2963, B => n9, C => n2962, D => n180, Z => n737)
                           ;
   U3309 : NR4 port map( A => n739, B => n740, C => n741, D => n742, Z => n733)
                           ;
   U3310 : AO4 port map( A => n2967, B => n53, C => n2966, D => n170, Z => n739
                           );
   U3311 : AO4 port map( A => n2969, B => n249, C => n2968, D => n250, Z => 
                           n740);
   U3312 : AO4 port map( A => n2971, B => n28, C => n2970, D => n14, Z => n741)
                           ;
   U3313 : NR4 port map( A => n743, B => n744, C => n745, D => n746, Z => n732)
                           ;
   U3314 : AO4 port map( A => n2975, B => n8, C => n2974, D => n163, Z => n743)
                           ;
   U3315 : AO4 port map( A => n2977, B => n258, C => n2976, D => n259, Z => 
                           n744);
   U3316 : AO4 port map( A => n2979, B => n7, C => n2978, D => n150, Z => n745)
                           ;
   U3317 : NR4 port map( A => n747, B => n748, C => n749, D => n750, Z => n731)
                           ;
   U3318 : AO4 port map( A => n2983, B => n48, C => n2982, D => n122, Z => n747
                           );
   U3319 : AO4 port map( A => n2985, B => n246, C => n2984, D => n248, Z => 
                           n748);
   U3320 : AO4 port map( A => n2987, B => n6, C => n2986, D => n109, Z => n749)
                           ;
   U3321 : NR4 port map( A => n759, B => n760, C => n761, D => n762, Z => n758)
                           ;
   U3322 : AO4 port map( A => n3055, B => n81, C => n3054, D => n229, Z => n759
                           );
   U3323 : AO4 port map( A => n3057, B => n270, C => n3056, D => n272, Z => 
                           n760);
   U3324 : AO4 port map( A => n3059, B => n72, C => n3058, D => n228, Z => n761
                           );
   U3325 : NR4 port map( A => n763, B => n764, C => n765, D => n766, Z => n757)
                           ;
   U3326 : AO4 port map( A => n3063, B => n71, C => n3062, D => n227, Z => n763
                           );
   U3327 : AO4 port map( A => n3065, B => n255, C => n3064, D => n257, Z => 
                           n764);
   U3328 : AO4 port map( A => n3067, B => n12, C => n3066, D => n23, Z => n765)
                           ;
   U3329 : NR4 port map( A => n767, B => n768, C => n769, D => n770, Z => n756)
                           ;
   U3330 : AO4 port map( A => n3071, B => n69, C => n3070, D => n224, Z => n767
                           );
   U3331 : AO4 port map( A => n3073, B => n265, C => n3072, D => n269, Z => 
                           n768);
   U3332 : AO4 port map( A => n3075, B => n11, C => n3074, D => n217, Z => n769
                           );
   U3333 : NR4 port map( A => n771, B => n772, C => n773, D => n774, Z => n755)
                           ;
   U3334 : AO4 port map( A => n3079, B => n59, C => n3078, D => n209, Z => n771
                           );
   U3335 : AO4 port map( A => n3081, B => n251, C => n3080, D => n253, Z => 
                           n772);
   U3336 : AO4 port map( A => n3083, B => n10, C => n3082, D => n22, Z => n773)
                           ;
   U3337 : NR4 port map( A => n779, B => n780, C => n781, D => n782, Z => n778)
                           ;
   U3338 : AO4 port map( A => n3023, B => n58, C => n3022, D => n200, Z => n779
                           );
   U3339 : AO4 port map( A => n3025, B => n260, C => n3024, D => n261, Z => 
                           n780);
   U3340 : AO4 port map( A => n3027, B => n9, C => n3026, D => n180, Z => n781)
                           ;
   U3341 : NR4 port map( A => n783, B => n784, C => n785, D => n786, Z => n777)
                           ;
   U3342 : AO4 port map( A => n3031, B => n53, C => n3030, D => n170, Z => n783
                           );
   U3343 : AO4 port map( A => n3033, B => n249, C => n3032, D => n250, Z => 
                           n784);
   U3344 : AO4 port map( A => n3035, B => n28, C => n3034, D => n14, Z => n785)
                           ;
   U3345 : NR4 port map( A => n787, B => n788, C => n789, D => n790, Z => n776)
                           ;
   U3346 : AO4 port map( A => n3039, B => n8, C => n3038, D => n163, Z => n787)
                           ;
   U3347 : AO4 port map( A => n3041, B => n258, C => n3040, D => n259, Z => 
                           n788);
   U3348 : AO4 port map( A => n3043, B => n7, C => n3042, D => n150, Z => n789)
                           ;
   U3349 : NR4 port map( A => n791, B => n792, C => n793, D => n794, Z => n775)
                           ;
   U3350 : AO4 port map( A => n3047, B => n48, C => n3046, D => n122, Z => n791
                           );
   U3351 : AO4 port map( A => n3049, B => n246, C => n3048, D => n248, Z => 
                           n792);
   U3352 : AO4 port map( A => n3051, B => n6, C => n3050, D => n109, Z => n793)
                           ;
   U3353 : NR4 port map( A => n803, B => n804, C => n805, D => n806, Z => n802)
                           ;
   U3354 : AO4 port map( A => n3119, B => n81, C => n3118, D => n229, Z => n803
                           );
   U3355 : AO4 port map( A => n3121, B => n270, C => n3120, D => n272, Z => 
                           n804);
   U3356 : AO4 port map( A => n3123, B => n72, C => n3122, D => n228, Z => n805
                           );
   U3357 : NR4 port map( A => n807, B => n808, C => n809, D => n810, Z => n801)
                           ;
   U3358 : AO4 port map( A => n3127, B => n71, C => n3126, D => n227, Z => n807
                           );
   U3359 : AO4 port map( A => n3129, B => n255, C => n3128, D => n257, Z => 
                           n808);
   U3360 : AO4 port map( A => n3131, B => n12, C => n3130, D => n23, Z => n809)
                           ;
   U3361 : NR4 port map( A => n811, B => n812, C => n813, D => n814, Z => n800)
                           ;
   U3362 : AO4 port map( A => n3135, B => n69, C => n3134, D => n224, Z => n811
                           );
   U3363 : AO4 port map( A => n3137, B => n265, C => n3136, D => n269, Z => 
                           n812);
   U3364 : AO4 port map( A => n3139, B => n11, C => n3138, D => n217, Z => n813
                           );
   U3365 : NR4 port map( A => n815, B => n816, C => n817, D => n818, Z => n799)
                           ;
   U3366 : AO4 port map( A => n3143, B => n59, C => n3142, D => n209, Z => n815
                           );
   U3367 : AO4 port map( A => n3145, B => n251, C => n3144, D => n253, Z => 
                           n816);
   U3368 : AO4 port map( A => n3147, B => n10, C => n3146, D => n22, Z => n817)
                           ;
   U3369 : NR4 port map( A => n823, B => n824, C => n825, D => n826, Z => n822)
                           ;
   U3370 : AO4 port map( A => n3087, B => n58, C => n3086, D => n200, Z => n823
                           );
   U3371 : AO4 port map( A => n3089, B => n260, C => n3088, D => n261, Z => 
                           n824);
   U3372 : AO4 port map( A => n3091, B => n9, C => n3090, D => n180, Z => n825)
                           ;
   U3373 : NR4 port map( A => n827, B => n828, C => n829, D => n830, Z => n821)
                           ;
   U3374 : AO4 port map( A => n3095, B => n53, C => n3094, D => n170, Z => n827
                           );
   U3375 : AO4 port map( A => n3097, B => n249, C => n3096, D => n250, Z => 
                           n828);
   U3376 : AO4 port map( A => n3099, B => n28, C => n3098, D => n14, Z => n829)
                           ;
   U3377 : NR4 port map( A => n831, B => n832, C => n833, D => n834, Z => n820)
                           ;
   U3378 : AO4 port map( A => n3103, B => n8, C => n3102, D => n163, Z => n831)
                           ;
   U3379 : AO4 port map( A => n3105, B => n258, C => n3104, D => n259, Z => 
                           n832);
   U3380 : AO4 port map( A => n3107, B => n7, C => n3106, D => n150, Z => n833)
                           ;
   U3381 : NR4 port map( A => n835, B => n836, C => n837, D => n838, Z => n819)
                           ;
   U3382 : AO4 port map( A => n3111, B => n48, C => n3110, D => n122, Z => n835
                           );
   U3383 : AO4 port map( A => n3113, B => n246, C => n3112, D => n248, Z => 
                           n836);
   U3384 : AO4 port map( A => n3115, B => n6, C => n3114, D => n109, Z => n837)
                           ;
   U3385 : NR4 port map( A => n847, B => n848, C => n849, D => n850, Z => n846)
                           ;
   U3386 : AO4 port map( A => n3183, B => n81, C => n3182, D => n229, Z => n847
                           );
   U3387 : AO4 port map( A => n3185, B => n270, C => n3184, D => n272, Z => 
                           n848);
   U3388 : AO4 port map( A => n3187, B => n72, C => n3186, D => n228, Z => n849
                           );
   U3389 : NR4 port map( A => n851, B => n852, C => n853, D => n854, Z => n845)
                           ;
   U3390 : AO4 port map( A => n3191, B => n71, C => n3190, D => n227, Z => n851
                           );
   U3391 : AO4 port map( A => n3193, B => n255, C => n3192, D => n257, Z => 
                           n852);
   U3392 : AO4 port map( A => n3195, B => n12, C => n3194, D => n23, Z => n853)
                           ;
   U3393 : NR4 port map( A => n855, B => n856, C => n857, D => n858, Z => n844)
                           ;
   U3394 : AO4 port map( A => n3199, B => n69, C => n3198, D => n224, Z => n855
                           );
   U3395 : AO4 port map( A => n3201, B => n265, C => n3200, D => n269, Z => 
                           n856);
   U3396 : AO4 port map( A => n3203, B => n11, C => n3202, D => n217, Z => n857
                           );
   U3397 : NR4 port map( A => n859, B => n860, C => n861, D => n862, Z => n843)
                           ;
   U3398 : AO4 port map( A => n3207, B => n59, C => n3206, D => n209, Z => n859
                           );
   U3399 : AO4 port map( A => n3209, B => n251, C => n3208, D => n253, Z => 
                           n860);
   U3400 : AO4 port map( A => n3211, B => n10, C => n3210, D => n22, Z => n861)
                           ;
   U3401 : NR4 port map( A => n867, B => n868, C => n869, D => n870, Z => n866)
                           ;
   U3402 : AO4 port map( A => n3151, B => n58, C => n3150, D => n200, Z => n867
                           );
   U3403 : AO4 port map( A => n3153, B => n260, C => n3152, D => n261, Z => 
                           n868);
   U3404 : AO4 port map( A => n3155, B => n9, C => n3154, D => n180, Z => n869)
                           ;
   U3405 : NR4 port map( A => n871, B => n872, C => n873, D => n874, Z => n865)
                           ;
   U3406 : AO4 port map( A => n3159, B => n53, C => n3158, D => n170, Z => n871
                           );
   U3407 : AO4 port map( A => n3161, B => n249, C => n3160, D => n250, Z => 
                           n872);
   U3408 : AO4 port map( A => n3163, B => n28, C => n3162, D => n14, Z => n873)
                           ;
   U3409 : NR4 port map( A => n875, B => n876, C => n877, D => n878, Z => n864)
                           ;
   U3410 : AO4 port map( A => n3167, B => n8, C => n3166, D => n163, Z => n875)
                           ;
   U3411 : AO4 port map( A => n3169, B => n258, C => n3168, D => n259, Z => 
                           n876);
   U3412 : AO4 port map( A => n3171, B => n7, C => n3170, D => n150, Z => n877)
                           ;
   U3413 : NR4 port map( A => n879, B => n880, C => n881, D => n882, Z => n863)
                           ;
   U3414 : AO4 port map( A => n3175, B => n48, C => n3174, D => n122, Z => n879
                           );
   U3415 : AO4 port map( A => n3177, B => n246, C => n3176, D => n248, Z => 
                           n880);
   U3416 : AO4 port map( A => n3179, B => n6, C => n3178, D => n109, Z => n881)
                           ;
   U3417 : NR4 port map( A => n891, B => n892, C => n893, D => n894, Z => n890)
                           ;
   U3418 : AO4 port map( A => n3247, B => n81, C => n3246, D => n229, Z => n891
                           );
   U3419 : AO4 port map( A => n3249, B => n270, C => n3248, D => n272, Z => 
                           n892);
   U3420 : AO4 port map( A => n3251, B => n72, C => n3250, D => n228, Z => n893
                           );
   U3421 : NR4 port map( A => n895, B => n896, C => n897, D => n898, Z => n889)
                           ;
   U3422 : AO4 port map( A => n3255, B => n71, C => n3254, D => n227, Z => n895
                           );
   U3423 : AO4 port map( A => n3257, B => n255, C => n3256, D => n257, Z => 
                           n896);
   U3424 : AO4 port map( A => n3259, B => n12, C => n3258, D => n23, Z => n897)
                           ;
   U3425 : NR4 port map( A => n899, B => n900, C => n901, D => n902, Z => n888)
                           ;
   U3426 : AO4 port map( A => n3263, B => n69, C => n3262, D => n224, Z => n899
                           );
   U3427 : AO4 port map( A => n3265, B => n265, C => n3264, D => n269, Z => 
                           n900);
   U3428 : AO4 port map( A => n3267, B => n11, C => n3266, D => n217, Z => n901
                           );
   U3429 : NR4 port map( A => n903, B => n904, C => n905, D => n906, Z => n887)
                           ;
   U3430 : AO4 port map( A => n3271, B => n59, C => n3270, D => n209, Z => n903
                           );
   U3431 : AO4 port map( A => n3273, B => n251, C => n3272, D => n253, Z => 
                           n904);
   U3432 : AO4 port map( A => n3275, B => n10, C => n3274, D => n22, Z => n905)
                           ;
   U3433 : NR4 port map( A => n911, B => n912, C => n913, D => n914, Z => n910)
                           ;
   U3434 : AO4 port map( A => n3215, B => n58, C => n3214, D => n200, Z => n911
                           );
   U3435 : AO4 port map( A => n3217, B => n260, C => n3216, D => n261, Z => 
                           n912);
   U3436 : AO4 port map( A => n3219, B => n9, C => n3218, D => n180, Z => n913)
                           ;
   U3437 : NR4 port map( A => n915, B => n916, C => n917, D => n918, Z => n909)
                           ;
   U3438 : AO4 port map( A => n3223, B => n53, C => n3222, D => n170, Z => n915
                           );
   U3439 : AO4 port map( A => n3225, B => n249, C => n3224, D => n250, Z => 
                           n916);
   U3440 : AO4 port map( A => n3227, B => n28, C => n3226, D => n14, Z => n917)
                           ;
   U3441 : NR4 port map( A => n919, B => n920, C => n921, D => n922, Z => n908)
                           ;
   U3442 : AO4 port map( A => n3231, B => n8, C => n3230, D => n163, Z => n919)
                           ;
   U3443 : AO4 port map( A => n3233, B => n258, C => n3232, D => n259, Z => 
                           n920);
   U3444 : AO4 port map( A => n3235, B => n7, C => n3234, D => n150, Z => n921)
                           ;
   U3445 : NR4 port map( A => n923, B => n924, C => n925, D => n926, Z => n907)
                           ;
   U3446 : AO4 port map( A => n3239, B => n48, C => n3238, D => n122, Z => n923
                           );
   U3447 : AO4 port map( A => n3241, B => n246, C => n3240, D => n248, Z => 
                           n924);
   U3448 : AO4 port map( A => n3243, B => n6, C => n3242, D => n109, Z => n925)
                           ;
   U3449 : NR4 port map( A => n935, B => n936, C => n937, D => n938, Z => n934)
                           ;
   U3450 : AO4 port map( A => n3311, B => n81, C => n3310, D => n229, Z => n935
                           );
   U3451 : AO4 port map( A => n3313, B => n270, C => n3312, D => n272, Z => 
                           n936);
   U3452 : AO4 port map( A => n3315, B => n72, C => n3314, D => n228, Z => n937
                           );
   U3453 : NR4 port map( A => n939, B => n940, C => n941, D => n942, Z => n933)
                           ;
   U3454 : AO4 port map( A => n3319, B => n71, C => n3318, D => n227, Z => n939
                           );
   U3455 : AO4 port map( A => n3321, B => n255, C => n3320, D => n257, Z => 
                           n940);
   U3456 : AO4 port map( A => n3323, B => n12, C => n3322, D => n23, Z => n941)
                           ;
   U3457 : NR4 port map( A => n943, B => n944, C => n945, D => n946, Z => n932)
                           ;
   U3458 : AO4 port map( A => n3327, B => n69, C => n3326, D => n224, Z => n943
                           );
   U3459 : AO4 port map( A => n3329, B => n265, C => n3328, D => n269, Z => 
                           n944);
   U3460 : AO4 port map( A => n3331, B => n11, C => n3330, D => n217, Z => n945
                           );
   U3461 : NR4 port map( A => n947, B => n948, C => n949, D => n950, Z => n931)
                           ;
   U3462 : AO4 port map( A => n3335, B => n59, C => n3334, D => n209, Z => n947
                           );
   U3463 : AO4 port map( A => n3337, B => n251, C => n3336, D => n253, Z => 
                           n948);
   U3464 : AO4 port map( A => n3339, B => n10, C => n3338, D => n22, Z => n949)
                           ;
   U3465 : NR4 port map( A => n955, B => n956, C => n957, D => n958, Z => n954)
                           ;
   U3466 : AO4 port map( A => n3279, B => n58, C => n3278, D => n200, Z => n955
                           );
   U3467 : AO4 port map( A => n3281, B => n260, C => n3280, D => n261, Z => 
                           n956);
   U3468 : AO4 port map( A => n3283, B => n9, C => n3282, D => n180, Z => n957)
                           ;
   U3469 : NR4 port map( A => n959, B => n960, C => n961, D => n962, Z => n953)
                           ;
   U3470 : AO4 port map( A => n3287, B => n53, C => n3286, D => n170, Z => n959
                           );
   U3471 : AO4 port map( A => n3289, B => n249, C => n3288, D => n250, Z => 
                           n960);
   U3472 : AO4 port map( A => n3291, B => n28, C => n3290, D => n14, Z => n961)
                           ;
   U3473 : NR4 port map( A => n963, B => n964, C => n965, D => n966, Z => n952)
                           ;
   U3474 : AO4 port map( A => n3295, B => n8, C => n3294, D => n163, Z => n963)
                           ;
   U3475 : AO4 port map( A => n3297, B => n258, C => n3296, D => n259, Z => 
                           n964);
   U3476 : AO4 port map( A => n3299, B => n7, C => n3298, D => n150, Z => n965)
                           ;
   U3477 : NR4 port map( A => n967, B => n968, C => n969, D => n970, Z => n951)
                           ;
   U3478 : AO4 port map( A => n3303, B => n48, C => n3302, D => n122, Z => n967
                           );
   U3479 : AO4 port map( A => n3305, B => n246, C => n3304, D => n248, Z => 
                           n968);
   U3480 : AO4 port map( A => n3307, B => n6, C => n3306, D => n109, Z => n969)
                           ;
   U3481 : NR4 port map( A => n979, B => n980, C => n981, D => n982, Z => n978)
                           ;
   U3482 : AO4 port map( A => n3375, B => n81, C => n3374, D => n229, Z => n979
                           );
   U3483 : AO4 port map( A => n3377, B => n270, C => n3376, D => n272, Z => 
                           n980);
   U3484 : AO4 port map( A => n3379, B => n72, C => n3378, D => n228, Z => n981
                           );
   U3485 : NR4 port map( A => n983, B => n984, C => n985, D => n986, Z => n977)
                           ;
   U3486 : AO4 port map( A => n3383, B => n71, C => n3382, D => n227, Z => n983
                           );
   U3487 : AO4 port map( A => n3385, B => n255, C => n3384, D => n257, Z => 
                           n984);
   U3488 : AO4 port map( A => n3387, B => n12, C => n3386, D => n23, Z => n985)
                           ;
   U3489 : NR4 port map( A => n987, B => n988, C => n989, D => n990, Z => n976)
                           ;
   U3490 : AO4 port map( A => n3391, B => n69, C => n3390, D => n224, Z => n987
                           );
   U3491 : AO4 port map( A => n3393, B => n265, C => n3392, D => n269, Z => 
                           n988);
   U3492 : AO4 port map( A => n3395, B => n11, C => n3394, D => n217, Z => n989
                           );
   U3493 : NR4 port map( A => n991, B => n992, C => n993, D => n994, Z => n975)
                           ;
   U3494 : AO4 port map( A => n3399, B => n59, C => n3398, D => n209, Z => n991
                           );
   U3495 : AO4 port map( A => n3401, B => n251, C => n3400, D => n253, Z => 
                           n992);
   U3496 : AO4 port map( A => n3403, B => n10, C => n3402, D => n22, Z => n993)
                           ;
   U3497 : NR4 port map( A => n999, B => n1000, C => n1001, D => n1002, Z => 
                           n998);
   U3498 : AO4 port map( A => n3343, B => n58, C => n3342, D => n200, Z => n999
                           );
   U3499 : AO4 port map( A => n3345, B => n260, C => n3344, D => n261, Z => 
                           n1000);
   U3500 : AO4 port map( A => n3347, B => n9, C => n3346, D => n180, Z => n1001
                           );
   U3501 : NR4 port map( A => n1003, B => n1004, C => n1005, D => n1006, Z => 
                           n997);
   U3502 : AO4 port map( A => n3351, B => n53, C => n3350, D => n170, Z => 
                           n1003);
   U3503 : AO4 port map( A => n3353, B => n249, C => n3352, D => n250, Z => 
                           n1004);
   U3504 : AO4 port map( A => n3355, B => n28, C => n3354, D => n14, Z => n1005
                           );
   U3505 : NR4 port map( A => n1007, B => n1008, C => n1009, D => n1010, Z => 
                           n996);
   U3506 : AO4 port map( A => n3359, B => n8, C => n3358, D => n163, Z => n1007
                           );
   U3507 : AO4 port map( A => n3361, B => n258, C => n3360, D => n259, Z => 
                           n1008);
   U3508 : AO4 port map( A => n3363, B => n7, C => n3362, D => n150, Z => n1009
                           );
   U3509 : NR4 port map( A => n1011, B => n1012, C => n1013, D => n1014, Z => 
                           n995);
   U3510 : AO4 port map( A => n3367, B => n48, C => n3366, D => n122, Z => 
                           n1011);
   U3511 : AO4 port map( A => n3369, B => n246, C => n3368, D => n248, Z => 
                           n1012);
   U3512 : AO4 port map( A => n3371, B => n6, C => n3370, D => n109, Z => n1013
                           );
   U3513 : NR4 port map( A => n1023, B => n1024, C => n1025, D => n1026, Z => 
                           n1022);
   U3514 : AO4 port map( A => n3439, B => n81, C => n3438, D => n229, Z => 
                           n1023);
   U3515 : AO4 port map( A => n3441, B => n270, C => n3440, D => n272, Z => 
                           n1024);
   U3516 : AO4 port map( A => n3443, B => n72, C => n3442, D => n228, Z => 
                           n1025);
   U3517 : NR4 port map( A => n1027, B => n1028, C => n1029, D => n1030, Z => 
                           n1021);
   U3518 : AO4 port map( A => n3447, B => n71, C => n3446, D => n227, Z => 
                           n1027);
   U3519 : AO4 port map( A => n3449, B => n255, C => n3448, D => n257, Z => 
                           n1028);
   U3520 : AO4 port map( A => n3451, B => n12, C => n3450, D => n23, Z => n1029
                           );
   U3521 : NR4 port map( A => n1031, B => n1032, C => n1033, D => n1034, Z => 
                           n1020);
   U3522 : AO4 port map( A => n3455, B => n69, C => n3454, D => n224, Z => 
                           n1031);
   U3523 : AO4 port map( A => n3457, B => n265, C => n3456, D => n269, Z => 
                           n1032);
   U3524 : AO4 port map( A => n3459, B => n11, C => n3458, D => n217, Z => 
                           n1033);
   U3525 : NR4 port map( A => n1035, B => n1036, C => n1037, D => n1038, Z => 
                           n1019);
   U3526 : AO4 port map( A => n3463, B => n59, C => n3462, D => n209, Z => 
                           n1035);
   U3527 : AO4 port map( A => n3465, B => n251, C => n3464, D => n253, Z => 
                           n1036);
   U3528 : AO4 port map( A => n3467, B => n10, C => n3466, D => n22, Z => n1037
                           );
   U3529 : NR4 port map( A => n1043, B => n1044, C => n1045, D => n1046, Z => 
                           n1042);
   U3530 : AO4 port map( A => n3407, B => n58, C => n3406, D => n200, Z => 
                           n1043);
   U3531 : AO4 port map( A => n3409, B => n260, C => n3408, D => n261, Z => 
                           n1044);
   U3532 : AO4 port map( A => n3411, B => n9, C => n3410, D => n180, Z => n1045
                           );
   U3533 : NR4 port map( A => n1047, B => n1048, C => n1049, D => n1050, Z => 
                           n1041);
   U3534 : AO4 port map( A => n3415, B => n53, C => n3414, D => n170, Z => 
                           n1047);
   U3535 : AO4 port map( A => n3417, B => n249, C => n3416, D => n250, Z => 
                           n1048);
   U3536 : AO4 port map( A => n3419, B => n28, C => n3418, D => n14, Z => n1049
                           );
   U3537 : NR4 port map( A => n1051, B => n1052, C => n1053, D => n1054, Z => 
                           n1040);
   U3538 : AO4 port map( A => n3423, B => n8, C => n3422, D => n163, Z => n1051
                           );
   U3539 : AO4 port map( A => n3425, B => n258, C => n3424, D => n259, Z => 
                           n1052);
   U3540 : AO4 port map( A => n3427, B => n7, C => n3426, D => n150, Z => n1053
                           );
   U3541 : NR4 port map( A => n1055, B => n1056, C => n1057, D => n1058, Z => 
                           n1039);
   U3542 : AO4 port map( A => n3431, B => n48, C => n3430, D => n122, Z => 
                           n1055);
   U3543 : AO4 port map( A => n3433, B => n246, C => n3432, D => n248, Z => 
                           n1056);
   U3544 : AO4 port map( A => n3435, B => n6, C => n3434, D => n109, Z => n1057
                           );
   U3545 : NR4 port map( A => n1067, B => n1068, C => n1069, D => n1070, Z => 
                           n1066);
   U3546 : AO4 port map( A => n3503, B => n81, C => n3502, D => n229, Z => 
                           n1067);
   U3547 : AO4 port map( A => n3505, B => n270, C => n3504, D => n272, Z => 
                           n1068);
   U3548 : AO4 port map( A => n3507, B => n72, C => n3506, D => n228, Z => 
                           n1069);
   U3549 : NR4 port map( A => n1071, B => n1072, C => n1073, D => n1074, Z => 
                           n1065);
   U3550 : AO4 port map( A => n3511, B => n71, C => n3510, D => n227, Z => 
                           n1071);
   U3551 : AO4 port map( A => n3513, B => n255, C => n3512, D => n257, Z => 
                           n1072);
   U3552 : AO4 port map( A => n3515, B => n12, C => n3514, D => n23, Z => n1073
                           );
   U3553 : NR4 port map( A => n1075, B => n1076, C => n1077, D => n1078, Z => 
                           n1064);
   U3554 : AO4 port map( A => n3519, B => n69, C => n3518, D => n224, Z => 
                           n1075);
   U3555 : AO4 port map( A => n3521, B => n265, C => n3520, D => n269, Z => 
                           n1076);
   U3556 : AO4 port map( A => n3523, B => n11, C => n3522, D => n217, Z => 
                           n1077);
   U3557 : NR4 port map( A => n1079, B => n1080, C => n1081, D => n1082, Z => 
                           n1063);
   U3558 : AO4 port map( A => n3527, B => n59, C => n3526, D => n209, Z => 
                           n1079);
   U3559 : AO4 port map( A => n3529, B => n251, C => n3528, D => n253, Z => 
                           n1080);
   U3560 : AO4 port map( A => n3531, B => n10, C => n3530, D => n22, Z => n1081
                           );
   U3561 : NR4 port map( A => n1087, B => n1088, C => n1089, D => n1090, Z => 
                           n1086);
   U3562 : AO4 port map( A => n3471, B => n58, C => n3470, D => n200, Z => 
                           n1087);
   U3563 : AO4 port map( A => n3473, B => n260, C => n3472, D => n261, Z => 
                           n1088);
   U3564 : AO4 port map( A => n3475, B => n9, C => n3474, D => n180, Z => n1089
                           );
   U3565 : NR4 port map( A => n1091, B => n1092, C => n1093, D => n1094, Z => 
                           n1085);
   U3566 : AO4 port map( A => n3479, B => n53, C => n3478, D => n170, Z => 
                           n1091);
   U3567 : AO4 port map( A => n3481, B => n249, C => n3480, D => n250, Z => 
                           n1092);
   U3568 : AO4 port map( A => n3483, B => n28, C => n3482, D => n14, Z => n1093
                           );
   U3569 : NR4 port map( A => n1095, B => n1096, C => n1097, D => n1098, Z => 
                           n1084);
   U3570 : AO4 port map( A => n3487, B => n8, C => n3486, D => n163, Z => n1095
                           );
   U3571 : AO4 port map( A => n3489, B => n258, C => n3488, D => n259, Z => 
                           n1096);
   U3572 : AO4 port map( A => n3491, B => n7, C => n3490, D => n150, Z => n1097
                           );
   U3573 : NR4 port map( A => n1099, B => n1100, C => n1101, D => n1102, Z => 
                           n1083);
   U3574 : AO4 port map( A => n3495, B => n48, C => n3494, D => n122, Z => 
                           n1099);
   U3575 : AO4 port map( A => n3497, B => n246, C => n3496, D => n248, Z => 
                           n1100);
   U3576 : AO4 port map( A => n3499, B => n6, C => n3498, D => n109, Z => n1101
                           );
   U3577 : NR4 port map( A => n1111, B => n1112, C => n1113, D => n1114, Z => 
                           n1110);
   U3578 : AO4 port map( A => n3567, B => n81, C => n3566, D => n229, Z => 
                           n1111);
   U3579 : AO4 port map( A => n3569, B => n270, C => n3568, D => n272, Z => 
                           n1112);
   U3580 : AO4 port map( A => n3571, B => n72, C => n3570, D => n228, Z => 
                           n1113);
   U3581 : NR4 port map( A => n1115, B => n1116, C => n1117, D => n1118, Z => 
                           n1109);
   U3582 : AO4 port map( A => n3575, B => n71, C => n3574, D => n227, Z => 
                           n1115);
   U3583 : AO4 port map( A => n3577, B => n255, C => n3576, D => n257, Z => 
                           n1116);
   U3584 : AO4 port map( A => n3579, B => n12, C => n3578, D => n23, Z => n1117
                           );
   U3585 : NR4 port map( A => n1119, B => n1120, C => n1121, D => n1122, Z => 
                           n1108);
   U3586 : AO4 port map( A => n3583, B => n69, C => n3582, D => n224, Z => 
                           n1119);
   U3587 : AO4 port map( A => n3585, B => n265, C => n3584, D => n269, Z => 
                           n1120);
   U3588 : AO4 port map( A => n3587, B => n11, C => n3586, D => n217, Z => 
                           n1121);
   U3589 : NR4 port map( A => n1123, B => n1124, C => n1125, D => n1126, Z => 
                           n1107);
   U3590 : AO4 port map( A => n3591, B => n59, C => n3590, D => n209, Z => 
                           n1123);
   U3591 : AO4 port map( A => n3593, B => n251, C => n3592, D => n253, Z => 
                           n1124);
   U3592 : AO4 port map( A => n3595, B => n10, C => n3594, D => n22, Z => n1125
                           );
   U3593 : NR4 port map( A => n1131, B => n1132, C => n1133, D => n1134, Z => 
                           n1130);
   U3594 : AO4 port map( A => n3535, B => n58, C => n3534, D => n200, Z => 
                           n1131);
   U3595 : AO4 port map( A => n3537, B => n260, C => n3536, D => n261, Z => 
                           n1132);
   U3596 : AO4 port map( A => n3539, B => n9, C => n3538, D => n180, Z => n1133
                           );
   U3597 : NR4 port map( A => n1135, B => n1136, C => n1137, D => n1138, Z => 
                           n1129);
   U3598 : AO4 port map( A => n3543, B => n53, C => n3542, D => n170, Z => 
                           n1135);
   U3599 : AO4 port map( A => n3545, B => n249, C => n3544, D => n250, Z => 
                           n1136);
   U3600 : AO4 port map( A => n3547, B => n28, C => n3546, D => n14, Z => n1137
                           );
   U3601 : NR4 port map( A => n1139, B => n1140, C => n1141, D => n1142, Z => 
                           n1128);
   U3602 : AO4 port map( A => n3551, B => n8, C => n3550, D => n163, Z => n1139
                           );
   U3603 : AO4 port map( A => n3553, B => n258, C => n3552, D => n259, Z => 
                           n1140);
   U3604 : AO4 port map( A => n3555, B => n7, C => n3554, D => n150, Z => n1141
                           );
   U3605 : NR4 port map( A => n1143, B => n1144, C => n1145, D => n1146, Z => 
                           n1127);
   U3606 : AO4 port map( A => n3559, B => n48, C => n3558, D => n122, Z => 
                           n1143);
   U3607 : AO4 port map( A => n3561, B => n246, C => n3560, D => n248, Z => 
                           n1144);
   U3608 : AO4 port map( A => n3563, B => n6, C => n3562, D => n109, Z => n1145
                           );
   U3609 : NR4 port map( A => n1155, B => n1156, C => n1157, D => n1158, Z => 
                           n1154);
   U3610 : AO4 port map( A => n3631, B => n81, C => n3630, D => n229, Z => 
                           n1155);
   U3611 : AO4 port map( A => n3633, B => n270, C => n3632, D => n272, Z => 
                           n1156);
   U3612 : AO4 port map( A => n3635, B => n72, C => n3634, D => n228, Z => 
                           n1157);
   U3613 : NR4 port map( A => n1159, B => n1160, C => n1161, D => n1162, Z => 
                           n1153);
   U3614 : AO4 port map( A => n3639, B => n71, C => n3638, D => n227, Z => 
                           n1159);
   U3615 : AO4 port map( A => n3641, B => n255, C => n3640, D => n257, Z => 
                           n1160);
   U3616 : AO4 port map( A => n3643, B => n12, C => n3642, D => n23, Z => n1161
                           );
   U3617 : NR4 port map( A => n1163, B => n1164, C => n1165, D => n1166, Z => 
                           n1152);
   U3618 : AO4 port map( A => n3647, B => n69, C => n3646, D => n224, Z => 
                           n1163);
   U3619 : AO4 port map( A => n3649, B => n265, C => n3648, D => n269, Z => 
                           n1164);
   U3620 : AO4 port map( A => n3651, B => n11, C => n3650, D => n217, Z => 
                           n1165);
   U3621 : NR4 port map( A => n1167, B => n1168, C => n1169, D => n1170, Z => 
                           n1151);
   U3622 : AO4 port map( A => n3655, B => n59, C => n3654, D => n209, Z => 
                           n1167);
   U3623 : AO4 port map( A => n3657, B => n251, C => n3656, D => n253, Z => 
                           n1168);
   U3624 : AO4 port map( A => n3659, B => n10, C => n3658, D => n22, Z => n1169
                           );
   U3625 : NR4 port map( A => n1175, B => n1176, C => n1177, D => n1178, Z => 
                           n1174);
   U3626 : AO4 port map( A => n3599, B => n58, C => n3598, D => n200, Z => 
                           n1175);
   U3627 : AO4 port map( A => n3601, B => n260, C => n3600, D => n261, Z => 
                           n1176);
   U3628 : AO4 port map( A => n3603, B => n9, C => n3602, D => n180, Z => n1177
                           );
   U3629 : NR4 port map( A => n1179, B => n1180, C => n1181, D => n1182, Z => 
                           n1173);
   U3630 : AO4 port map( A => n3607, B => n53, C => n3606, D => n170, Z => 
                           n1179);
   U3631 : AO4 port map( A => n3609, B => n249, C => n3608, D => n250, Z => 
                           n1180);
   U3632 : AO4 port map( A => n3611, B => n28, C => n3610, D => n14, Z => n1181
                           );
   U3633 : NR4 port map( A => n1183, B => n1184, C => n1185, D => n1186, Z => 
                           n1172);
   U3634 : AO4 port map( A => n3615, B => n8, C => n3614, D => n163, Z => n1183
                           );
   U3635 : AO4 port map( A => n3617, B => n258, C => n3616, D => n259, Z => 
                           n1184);
   U3636 : AO4 port map( A => n3619, B => n7, C => n3618, D => n150, Z => n1185
                           );
   U3637 : NR4 port map( A => n1187, B => n1188, C => n1189, D => n1190, Z => 
                           n1171);
   U3638 : AO4 port map( A => n3623, B => n48, C => n3622, D => n122, Z => 
                           n1187);
   U3639 : AO4 port map( A => n3625, B => n246, C => n3624, D => n248, Z => 
                           n1188);
   U3640 : AO4 port map( A => n3627, B => n6, C => n3626, D => n109, Z => n1189
                           );
   U3641 : NR4 port map( A => n1199, B => n1200, C => n1201, D => n1202, Z => 
                           n1198);
   U3642 : AO4 port map( A => n3695, B => n81, C => n3694, D => n229, Z => 
                           n1199);
   U3643 : AO4 port map( A => n3697, B => n270, C => n3696, D => n272, Z => 
                           n1200);
   U3644 : AO4 port map( A => n3699, B => n72, C => n3698, D => n228, Z => 
                           n1201);
   U3645 : NR4 port map( A => n1203, B => n1204, C => n1205, D => n1206, Z => 
                           n1197);
   U3646 : AO4 port map( A => n3703, B => n71, C => n3702, D => n227, Z => 
                           n1203);
   U3647 : AO4 port map( A => n3705, B => n255, C => n3704, D => n257, Z => 
                           n1204);
   U3648 : AO4 port map( A => n3707, B => n12, C => n3706, D => n23, Z => n1205
                           );
   U3649 : NR4 port map( A => n1207, B => n1208, C => n1209, D => n1210, Z => 
                           n1196);
   U3650 : AO4 port map( A => n3711, B => n69, C => n3710, D => n224, Z => 
                           n1207);
   U3651 : AO4 port map( A => n3713, B => n265, C => n3712, D => n269, Z => 
                           n1208);
   U3652 : AO4 port map( A => n3715, B => n11, C => n3714, D => n217, Z => 
                           n1209);
   U3653 : NR4 port map( A => n1211, B => n1212, C => n1213, D => n1214, Z => 
                           n1195);
   U3654 : AO4 port map( A => n3719, B => n59, C => n3718, D => n209, Z => 
                           n1211);
   U3655 : AO4 port map( A => n3721, B => n251, C => n3720, D => n253, Z => 
                           n1212);
   U3656 : AO4 port map( A => n3723, B => n10, C => n3722, D => n22, Z => n1213
                           );
   U3657 : NR4 port map( A => n1219, B => n1220, C => n1221, D => n1222, Z => 
                           n1218);
   U3658 : AO4 port map( A => n3663, B => n58, C => n3662, D => n200, Z => 
                           n1219);
   U3659 : AO4 port map( A => n3665, B => n260, C => n3664, D => n261, Z => 
                           n1220);
   U3660 : AO4 port map( A => n3667, B => n9, C => n3666, D => n180, Z => n1221
                           );
   U3661 : NR4 port map( A => n1223, B => n1224, C => n1225, D => n1226, Z => 
                           n1217);
   U3662 : AO4 port map( A => n3671, B => n53, C => n3670, D => n170, Z => 
                           n1223);
   U3663 : AO4 port map( A => n3673, B => n249, C => n3672, D => n250, Z => 
                           n1224);
   U3664 : AO4 port map( A => n3675, B => n28, C => n3674, D => n14, Z => n1225
                           );
   U3665 : NR4 port map( A => n1227, B => n1228, C => n1229, D => n1230, Z => 
                           n1216);
   U3666 : AO4 port map( A => n3679, B => n8, C => n3678, D => n163, Z => n1227
                           );
   U3667 : AO4 port map( A => n3681, B => n258, C => n3680, D => n259, Z => 
                           n1228);
   U3668 : AO4 port map( A => n3683, B => n7, C => n3682, D => n150, Z => n1229
                           );
   U3669 : NR4 port map( A => n1231, B => n1232, C => n1233, D => n1234, Z => 
                           n1215);
   U3670 : AO4 port map( A => n3687, B => n48, C => n3686, D => n122, Z => 
                           n1231);
   U3671 : AO4 port map( A => n3689, B => n246, C => n3688, D => n248, Z => 
                           n1232);
   U3672 : AO4 port map( A => n3691, B => n6, C => n3690, D => n109, Z => n1233
                           );
   U3673 : NR4 port map( A => n1243, B => n1244, C => n1245, D => n1246, Z => 
                           n1242);
   U3674 : AO4 port map( A => n3759, B => n81, C => n3758, D => n229, Z => 
                           n1243);
   U3675 : AO4 port map( A => n3761, B => n270, C => n3760, D => n272, Z => 
                           n1244);
   U3676 : AO4 port map( A => n3763, B => n72, C => n3762, D => n228, Z => 
                           n1245);
   U3677 : NR4 port map( A => n1247, B => n1248, C => n1249, D => n1250, Z => 
                           n1241);
   U3678 : AO4 port map( A => n3767, B => n71, C => n3766, D => n227, Z => 
                           n1247);
   U3679 : AO4 port map( A => n3769, B => n255, C => n3768, D => n257, Z => 
                           n1248);
   U3680 : AO4 port map( A => n3771, B => n12, C => n3770, D => n23, Z => n1249
                           );
   U3681 : NR4 port map( A => n1251, B => n1252, C => n1253, D => n1254, Z => 
                           n1240);
   U3682 : AO4 port map( A => n3775, B => n69, C => n3774, D => n224, Z => 
                           n1251);
   U3683 : AO4 port map( A => n3777, B => n265, C => n3776, D => n269, Z => 
                           n1252);
   U3684 : AO4 port map( A => n3779, B => n11, C => n3778, D => n217, Z => 
                           n1253);
   U3685 : NR4 port map( A => n1255, B => n1256, C => n1257, D => n1258, Z => 
                           n1239);
   U3686 : AO4 port map( A => n3783, B => n59, C => n3782, D => n209, Z => 
                           n1255);
   U3687 : AO4 port map( A => n3785, B => n251, C => n3784, D => n253, Z => 
                           n1256);
   U3688 : AO4 port map( A => n3787, B => n10, C => n3786, D => n22, Z => n1257
                           );
   U3689 : NR4 port map( A => n1263, B => n1264, C => n1265, D => n1266, Z => 
                           n1262);
   U3690 : AO4 port map( A => n3727, B => n58, C => n3726, D => n200, Z => 
                           n1263);
   U3691 : AO4 port map( A => n3729, B => n260, C => n3728, D => n261, Z => 
                           n1264);
   U3692 : AO4 port map( A => n3731, B => n9, C => n3730, D => n180, Z => n1265
                           );
   U3693 : NR4 port map( A => n1267, B => n1268, C => n1269, D => n1270, Z => 
                           n1261);
   U3694 : AO4 port map( A => n3735, B => n53, C => n3734, D => n170, Z => 
                           n1267);
   U3695 : AO4 port map( A => n3737, B => n249, C => n3736, D => n250, Z => 
                           n1268);
   U3696 : AO4 port map( A => n3739, B => n28, C => n3738, D => n14, Z => n1269
                           );
   U3697 : NR4 port map( A => n1271, B => n1272, C => n1273, D => n1274, Z => 
                           n1260);
   U3698 : AO4 port map( A => n3743, B => n8, C => n3742, D => n163, Z => n1271
                           );
   U3699 : AO4 port map( A => n3745, B => n258, C => n3744, D => n259, Z => 
                           n1272);
   U3700 : AO4 port map( A => n3747, B => n7, C => n3746, D => n150, Z => n1273
                           );
   U3701 : NR4 port map( A => n1275, B => n1276, C => n1277, D => n1278, Z => 
                           n1259);
   U3702 : AO4 port map( A => n3751, B => n48, C => n3750, D => n122, Z => 
                           n1275);
   U3703 : AO4 port map( A => n3753, B => n246, C => n3752, D => n248, Z => 
                           n1276);
   U3704 : AO4 port map( A => n3755, B => n6, C => n3754, D => n109, Z => n1277
                           );
   U3705 : NR4 port map( A => n1287, B => n1288, C => n1289, D => n1290, Z => 
                           n1286);
   U3706 : AO4 port map( A => n3823, B => n81, C => n3822, D => n229, Z => 
                           n1287);
   U3707 : AO4 port map( A => n3825, B => n270, C => n3824, D => n272, Z => 
                           n1288);
   U3708 : AO4 port map( A => n3827, B => n72, C => n3826, D => n228, Z => 
                           n1289);
   U3709 : NR4 port map( A => n1291, B => n1292, C => n1293, D => n1294, Z => 
                           n1285);
   U3710 : AO4 port map( A => n3831, B => n71, C => n3830, D => n227, Z => 
                           n1291);
   U3711 : AO4 port map( A => n3833, B => n255, C => n3832, D => n257, Z => 
                           n1292);
   U3712 : AO4 port map( A => n3835, B => n12, C => n3834, D => n23, Z => n1293
                           );
   U3713 : NR4 port map( A => n1295, B => n1296, C => n1297, D => n1298, Z => 
                           n1284);
   U3714 : AO4 port map( A => n3839, B => n69, C => n3838, D => n224, Z => 
                           n1295);
   U3715 : AO4 port map( A => n3841, B => n265, C => n3840, D => n269, Z => 
                           n1296);
   U3716 : AO4 port map( A => n3843, B => n11, C => n3842, D => n217, Z => 
                           n1297);
   U3717 : NR4 port map( A => n1299, B => n1300, C => n1301, D => n1302, Z => 
                           n1283);
   U3718 : AO4 port map( A => n3847, B => n59, C => n3846, D => n209, Z => 
                           n1299);
   U3719 : AO4 port map( A => n3849, B => n251, C => n3848, D => n253, Z => 
                           n1300);
   U3720 : AO4 port map( A => n3851, B => n10, C => n3850, D => n22, Z => n1301
                           );
   U3721 : NR4 port map( A => n1307, B => n1308, C => n1309, D => n1310, Z => 
                           n1306);
   U3722 : AO4 port map( A => n3791, B => n58, C => n3790, D => n200, Z => 
                           n1307);
   U3723 : AO4 port map( A => n3793, B => n260, C => n3792, D => n261, Z => 
                           n1308);
   U3724 : AO4 port map( A => n3795, B => n9, C => n3794, D => n180, Z => n1309
                           );
   U3725 : NR4 port map( A => n1311, B => n1312, C => n1313, D => n1314, Z => 
                           n1305);
   U3726 : AO4 port map( A => n3799, B => n53, C => n3798, D => n170, Z => 
                           n1311);
   U3727 : AO4 port map( A => n3801, B => n249, C => n3800, D => n250, Z => 
                           n1312);
   U3728 : AO4 port map( A => n3803, B => n28, C => n3802, D => n14, Z => n1313
                           );
   U3729 : NR4 port map( A => n1315, B => n1316, C => n1317, D => n1318, Z => 
                           n1304);
   U3730 : AO4 port map( A => n3807, B => n8, C => n3806, D => n163, Z => n1315
                           );
   U3731 : AO4 port map( A => n3809, B => n258, C => n3808, D => n259, Z => 
                           n1316);
   U3732 : AO4 port map( A => n3811, B => n7, C => n3810, D => n150, Z => n1317
                           );
   U3733 : NR4 port map( A => n1319, B => n1320, C => n1321, D => n1322, Z => 
                           n1303);
   U3734 : AO4 port map( A => n3815, B => n48, C => n3814, D => n122, Z => 
                           n1319);
   U3735 : AO4 port map( A => n3817, B => n246, C => n3816, D => n248, Z => 
                           n1320);
   U3736 : AO4 port map( A => n3819, B => n6, C => n3818, D => n109, Z => n1321
                           );
   U3737 : NR4 port map( A => n1331, B => n1332, C => n1333, D => n1334, Z => 
                           n1330);
   U3738 : AO4 port map( A => n3887, B => n81, C => n3886, D => n229, Z => 
                           n1331);
   U3739 : AO4 port map( A => n3889, B => n270, C => n3888, D => n272, Z => 
                           n1332);
   U3740 : AO4 port map( A => n3891, B => n72, C => n3890, D => n228, Z => 
                           n1333);
   U3741 : NR4 port map( A => n1335, B => n1336, C => n1337, D => n1338, Z => 
                           n1329);
   U3742 : AO4 port map( A => n3895, B => n71, C => n3894, D => n227, Z => 
                           n1335);
   U3743 : AO4 port map( A => n3897, B => n255, C => n3896, D => n257, Z => 
                           n1336);
   U3744 : AO4 port map( A => n3899, B => n12, C => n3898, D => n23, Z => n1337
                           );
   U3745 : NR4 port map( A => n1339, B => n1340, C => n1341, D => n1342, Z => 
                           n1328);
   U3746 : AO4 port map( A => n3903, B => n69, C => n3902, D => n224, Z => 
                           n1339);
   U3747 : AO4 port map( A => n3905, B => n265, C => n3904, D => n269, Z => 
                           n1340);
   U3748 : AO4 port map( A => n3907, B => n11, C => n3906, D => n217, Z => 
                           n1341);
   U3749 : NR4 port map( A => n1343, B => n1344, C => n1345, D => n1346, Z => 
                           n1327);
   U3750 : AO4 port map( A => n3911, B => n59, C => n3910, D => n209, Z => 
                           n1343);
   U3751 : AO4 port map( A => n3913, B => n251, C => n3912, D => n253, Z => 
                           n1344);
   U3752 : AO4 port map( A => n3915, B => n10, C => n3914, D => n22, Z => n1345
                           );
   U3753 : NR4 port map( A => n1351, B => n1352, C => n1353, D => n1354, Z => 
                           n1350);
   U3754 : AO4 port map( A => n3855, B => n58, C => n3854, D => n200, Z => 
                           n1351);
   U3755 : AO4 port map( A => n3857, B => n260, C => n3856, D => n261, Z => 
                           n1352);
   U3756 : AO4 port map( A => n3859, B => n9, C => n3858, D => n180, Z => n1353
                           );
   U3757 : NR4 port map( A => n1355, B => n1356, C => n1357, D => n1358, Z => 
                           n1349);
   U3758 : AO4 port map( A => n3863, B => n53, C => n3862, D => n170, Z => 
                           n1355);
   U3759 : AO4 port map( A => n3865, B => n249, C => n3864, D => n250, Z => 
                           n1356);
   U3760 : AO4 port map( A => n3867, B => n28, C => n3866, D => n14, Z => n1357
                           );
   U3761 : NR4 port map( A => n1359, B => n1360, C => n1361, D => n1362, Z => 
                           n1348);
   U3762 : AO4 port map( A => n3871, B => n8, C => n3870, D => n163, Z => n1359
                           );
   U3763 : AO4 port map( A => n3873, B => n258, C => n3872, D => n259, Z => 
                           n1360);
   U3764 : AO4 port map( A => n3875, B => n7, C => n3874, D => n150, Z => n1361
                           );
   U3765 : NR4 port map( A => n1363, B => n1364, C => n1365, D => n1366, Z => 
                           n1347);
   U3766 : AO4 port map( A => n3879, B => n48, C => n3878, D => n122, Z => 
                           n1363);
   U3767 : AO4 port map( A => n3881, B => n246, C => n3880, D => n248, Z => 
                           n1364);
   U3768 : AO4 port map( A => n3883, B => n6, C => n3882, D => n109, Z => n1365
                           );
   U3769 : NR4 port map( A => n1375, B => n1376, C => n1377, D => n1378, Z => 
                           n1374);
   U3770 : AO4 port map( A => n3951, B => n81, C => n3950, D => n229, Z => 
                           n1375);
   U3771 : AO4 port map( A => n3953, B => n270, C => n3952, D => n272, Z => 
                           n1376);
   U3772 : AO4 port map( A => n3955, B => n72, C => n3954, D => n228, Z => 
                           n1377);
   U3773 : NR4 port map( A => n1379, B => n1380, C => n1381, D => n1382, Z => 
                           n1373);
   U3774 : AO4 port map( A => n3959, B => n71, C => n3958, D => n227, Z => 
                           n1379);
   U3775 : AO4 port map( A => n3961, B => n255, C => n3960, D => n257, Z => 
                           n1380);
   U3776 : AO4 port map( A => n3963, B => n12, C => n3962, D => n23, Z => n1381
                           );
   U3777 : NR4 port map( A => n1383, B => n1384, C => n1385, D => n1386, Z => 
                           n1372);
   U3778 : AO4 port map( A => n3967, B => n69, C => n3966, D => n224, Z => 
                           n1383);
   U3779 : AO4 port map( A => n3969, B => n265, C => n3968, D => n269, Z => 
                           n1384);
   U3780 : AO4 port map( A => n3971, B => n11, C => n3970, D => n217, Z => 
                           n1385);
   U3781 : NR4 port map( A => n1387, B => n1388, C => n1389, D => n1390, Z => 
                           n1371);
   U3782 : AO4 port map( A => n3975, B => n59, C => n3974, D => n209, Z => 
                           n1387);
   U3783 : AO4 port map( A => n3977, B => n251, C => n3976, D => n253, Z => 
                           n1388);
   U3784 : AO4 port map( A => n3979, B => n10, C => n3978, D => n22, Z => n1389
                           );
   U3785 : NR4 port map( A => n1395, B => n1396, C => n1397, D => n1398, Z => 
                           n1394);
   U3786 : AO4 port map( A => n3919, B => n58, C => n3918, D => n200, Z => 
                           n1395);
   U3787 : AO4 port map( A => n3921, B => n260, C => n3920, D => n261, Z => 
                           n1396);
   U3788 : AO4 port map( A => n3923, B => n9, C => n3922, D => n180, Z => n1397
                           );
   U3789 : NR4 port map( A => n1399, B => n1400, C => n1401, D => n1402, Z => 
                           n1393);
   U3790 : AO4 port map( A => n3927, B => n53, C => n3926, D => n170, Z => 
                           n1399);
   U3791 : AO4 port map( A => n3929, B => n249, C => n3928, D => n250, Z => 
                           n1400);
   U3792 : AO4 port map( A => n3931, B => n28, C => n3930, D => n14, Z => n1401
                           );
   U3793 : NR4 port map( A => n1403, B => n1404, C => n1405, D => n1406, Z => 
                           n1392);
   U3794 : AO4 port map( A => n3935, B => n8, C => n3934, D => n163, Z => n1403
                           );
   U3795 : AO4 port map( A => n3937, B => n258, C => n3936, D => n259, Z => 
                           n1404);
   U3796 : AO4 port map( A => n3939, B => n7, C => n3938, D => n150, Z => n1405
                           );
   U3797 : NR4 port map( A => n1407, B => n1408, C => n1409, D => n1410, Z => 
                           n1391);
   U3798 : AO4 port map( A => n3943, B => n48, C => n3942, D => n122, Z => 
                           n1407);
   U3799 : AO4 port map( A => n3945, B => n246, C => n3944, D => n248, Z => 
                           n1408);
   U3800 : AO4 port map( A => n3947, B => n6, C => n3946, D => n109, Z => n1409
                           );
   U3801 : NR4 port map( A => n1419, B => n1420, C => n1421, D => n1422, Z => 
                           n1418);
   U3802 : AO4 port map( A => n4015, B => n81, C => n4014, D => n229, Z => 
                           n1419);
   U3803 : AO4 port map( A => n4017, B => n270, C => n4016, D => n272, Z => 
                           n1420);
   U3804 : AO4 port map( A => n4019, B => n72, C => n4018, D => n228, Z => 
                           n1421);
   U3805 : NR4 port map( A => n1423, B => n1424, C => n1425, D => n1426, Z => 
                           n1417);
   U3806 : AO4 port map( A => n4023, B => n71, C => n4022, D => n227, Z => 
                           n1423);
   U3807 : AO4 port map( A => n4025, B => n255, C => n4024, D => n257, Z => 
                           n1424);
   U3808 : AO4 port map( A => n4027, B => n12, C => n4026, D => n23, Z => n1425
                           );
   U3809 : NR4 port map( A => n1427, B => n1428, C => n1429, D => n1430, Z => 
                           n1416);
   U3810 : AO4 port map( A => n4031, B => n69, C => n4030, D => n224, Z => 
                           n1427);
   U3811 : AO4 port map( A => n4033, B => n265, C => n4032, D => n269, Z => 
                           n1428);
   U3812 : AO4 port map( A => n4035, B => n11, C => n4034, D => n217, Z => 
                           n1429);
   U3813 : NR4 port map( A => n1431, B => n1432, C => n1433, D => n1434, Z => 
                           n1415);
   U3814 : AO4 port map( A => n4039, B => n59, C => n4038, D => n209, Z => 
                           n1431);
   U3815 : AO4 port map( A => n4041, B => n251, C => n4040, D => n253, Z => 
                           n1432);
   U3816 : AO4 port map( A => n4043, B => n10, C => n4042, D => n22, Z => n1433
                           );
   U3817 : NR4 port map( A => n1439, B => n1440, C => n1441, D => n1442, Z => 
                           n1438);
   U3818 : AO4 port map( A => n3983, B => n58, C => n3982, D => n200, Z => 
                           n1439);
   U3819 : AO4 port map( A => n3985, B => n260, C => n3984, D => n261, Z => 
                           n1440);
   U3820 : AO4 port map( A => n3987, B => n9, C => n3986, D => n180, Z => n1441
                           );
   U3821 : NR4 port map( A => n1443, B => n1444, C => n1445, D => n1446, Z => 
                           n1437);
   U3822 : AO4 port map( A => n3991, B => n53, C => n3990, D => n170, Z => 
                           n1443);
   U3823 : AO4 port map( A => n3993, B => n249, C => n3992, D => n250, Z => 
                           n1444);
   U3824 : AO4 port map( A => n3995, B => n28, C => n3994, D => n14, Z => n1445
                           );
   U3825 : NR4 port map( A => n1447, B => n1448, C => n1449, D => n1450, Z => 
                           n1436);
   U3826 : AO4 port map( A => n3999, B => n8, C => n3998, D => n163, Z => n1447
                           );
   U3827 : AO4 port map( A => n4001, B => n258, C => n4000, D => n259, Z => 
                           n1448);
   U3828 : AO4 port map( A => n4003, B => n7, C => n4002, D => n150, Z => n1449
                           );
   U3829 : NR4 port map( A => n1451, B => n1452, C => n1453, D => n1454, Z => 
                           n1435);
   U3830 : AO4 port map( A => n4007, B => n48, C => n4006, D => n122, Z => 
                           n1451);
   U3831 : AO4 port map( A => n4009, B => n246, C => n4008, D => n248, Z => 
                           n1452);
   U3832 : AO4 port map( A => n4011, B => n6, C => n4010, D => n109, Z => n1453
                           );
   U3833 : NR4 port map( A => n1463, B => n1464, C => n1465, D => n1466, Z => 
                           n1462);
   U3834 : AO4 port map( A => n4079, B => n81, C => n4078, D => n229, Z => 
                           n1463);
   U3835 : AO4 port map( A => n4081, B => n270, C => n4080, D => n272, Z => 
                           n1464);
   U3836 : AO4 port map( A => n4083, B => n72, C => n4082, D => n228, Z => 
                           n1465);
   U3837 : NR4 port map( A => n1467, B => n1468, C => n1469, D => n1470, Z => 
                           n1461);
   U3838 : AO4 port map( A => n4087, B => n71, C => n4086, D => n227, Z => 
                           n1467);
   U3839 : AO4 port map( A => n4089, B => n255, C => n4088, D => n257, Z => 
                           n1468);
   U3840 : AO4 port map( A => n4091, B => n12, C => n4090, D => n23, Z => n1469
                           );
   U3841 : NR4 port map( A => n1471, B => n1472, C => n1473, D => n1474, Z => 
                           n1460);
   U3842 : AO4 port map( A => n4095, B => n69, C => n4094, D => n224, Z => 
                           n1471);
   U3843 : AO4 port map( A => n4097, B => n265, C => n4096, D => n269, Z => 
                           n1472);
   U3844 : AO4 port map( A => n4099, B => n11, C => n4098, D => n217, Z => 
                           n1473);
   U3845 : NR4 port map( A => n1475, B => n1476, C => n1477, D => n1478, Z => 
                           n1459);
   U3846 : AO4 port map( A => n4103, B => n59, C => n4102, D => n209, Z => 
                           n1475);
   U3847 : AO4 port map( A => n4105, B => n251, C => n4104, D => n253, Z => 
                           n1476);
   U3848 : AO4 port map( A => n4107, B => n10, C => n4106, D => n22, Z => n1477
                           );
   U3849 : NR4 port map( A => n1483, B => n1484, C => n1485, D => n1486, Z => 
                           n1482);
   U3850 : AO4 port map( A => n4047, B => n58, C => n4046, D => n200, Z => 
                           n1483);
   U3851 : AO4 port map( A => n4049, B => n260, C => n4048, D => n261, Z => 
                           n1484);
   U3852 : AO4 port map( A => n4051, B => n9, C => n4050, D => n180, Z => n1485
                           );
   U3853 : NR4 port map( A => n1487, B => n1488, C => n1489, D => n1490, Z => 
                           n1481);
   U3854 : AO4 port map( A => n4055, B => n53, C => n4054, D => n170, Z => 
                           n1487);
   U3855 : AO4 port map( A => n4057, B => n249, C => n4056, D => n250, Z => 
                           n1488);
   U3856 : AO4 port map( A => n4059, B => n28, C => n4058, D => n14, Z => n1489
                           );
   U3857 : NR4 port map( A => n1491, B => n1492, C => n1493, D => n1494, Z => 
                           n1480);
   U3858 : AO4 port map( A => n4063, B => n8, C => n4062, D => n163, Z => n1491
                           );
   U3859 : AO4 port map( A => n4065, B => n258, C => n4064, D => n259, Z => 
                           n1492);
   U3860 : AO4 port map( A => n4067, B => n7, C => n4066, D => n150, Z => n1493
                           );
   U3861 : NR4 port map( A => n1495, B => n1496, C => n1497, D => n1498, Z => 
                           n1479);
   U3862 : AO4 port map( A => n4071, B => n48, C => n4070, D => n122, Z => 
                           n1495);
   U3863 : AO4 port map( A => n4073, B => n246, C => n4072, D => n248, Z => 
                           n1496);
   U3864 : AO4 port map( A => n4075, B => n6, C => n4074, D => n109, Z => n1497
                           );
   U3865 : NR4 port map( A => n1507, B => n1508, C => n1509, D => n1510, Z => 
                           n1506);
   U3866 : AO4 port map( A => n4143, B => n81, C => n4142, D => n229, Z => 
                           n1507);
   U3867 : AO4 port map( A => n4145, B => n270, C => n4144, D => n272, Z => 
                           n1508);
   U3868 : AO4 port map( A => n4147, B => n72, C => n4146, D => n228, Z => 
                           n1509);
   U3869 : NR4 port map( A => n1511, B => n1512, C => n1513, D => n1514, Z => 
                           n1505);
   U3870 : AO4 port map( A => n4151, B => n71, C => n4150, D => n227, Z => 
                           n1511);
   U3871 : AO4 port map( A => n4153, B => n255, C => n4152, D => n257, Z => 
                           n1512);
   U3872 : AO4 port map( A => n4155, B => n12, C => n4154, D => n23, Z => n1513
                           );
   U3873 : NR4 port map( A => n1515, B => n1516, C => n1517, D => n1518, Z => 
                           n1504);
   U3874 : AO4 port map( A => n4159, B => n69, C => n4158, D => n224, Z => 
                           n1515);
   U3875 : AO4 port map( A => n4161, B => n265, C => n4160, D => n269, Z => 
                           n1516);
   U3876 : AO4 port map( A => n4163, B => n11, C => n4162, D => n217, Z => 
                           n1517);
   U3877 : NR4 port map( A => n1519, B => n1520, C => n1521, D => n1522, Z => 
                           n1503);
   U3878 : AO4 port map( A => n4167, B => n59, C => n4166, D => n209, Z => 
                           n1519);
   U3879 : AO4 port map( A => n4169, B => n251, C => n4168, D => n253, Z => 
                           n1520);
   U3880 : AO4 port map( A => n4171, B => n10, C => n4170, D => n22, Z => n1521
                           );
   U3881 : NR4 port map( A => n1527, B => n1528, C => n1529, D => n1530, Z => 
                           n1526);
   U3882 : AO4 port map( A => n4111, B => n58, C => n4110, D => n200, Z => 
                           n1527);
   U3883 : AO4 port map( A => n4113, B => n260, C => n4112, D => n261, Z => 
                           n1528);
   U3884 : AO4 port map( A => n4115, B => n9, C => n4114, D => n180, Z => n1529
                           );
   U3885 : NR4 port map( A => n1531, B => n1532, C => n1533, D => n1534, Z => 
                           n1525);
   U3886 : AO4 port map( A => n4119, B => n53, C => n4118, D => n170, Z => 
                           n1531);
   U3887 : AO4 port map( A => n4121, B => n249, C => n4120, D => n250, Z => 
                           n1532);
   U3888 : AO4 port map( A => n4123, B => n28, C => n4122, D => n14, Z => n1533
                           );
   U3889 : NR4 port map( A => n1535, B => n1536, C => n1537, D => n1538, Z => 
                           n1524);
   U3890 : AO4 port map( A => n4127, B => n8, C => n4126, D => n163, Z => n1535
                           );
   U3891 : AO4 port map( A => n4129, B => n258, C => n4128, D => n259, Z => 
                           n1536);
   U3892 : AO4 port map( A => n4131, B => n7, C => n4130, D => n150, Z => n1537
                           );
   U3893 : NR4 port map( A => n1539, B => n1540, C => n1541, D => n1542, Z => 
                           n1523);
   U3894 : AO4 port map( A => n4135, B => n48, C => n4134, D => n122, Z => 
                           n1539);
   U3895 : AO4 port map( A => n4137, B => n246, C => n4136, D => n248, Z => 
                           n1540);
   U3896 : AO4 port map( A => n4139, B => n6, C => n4138, D => n109, Z => n1541
                           );
   U3897 : NR4 port map( A => n1551, B => n1552, C => n1553, D => n1554, Z => 
                           n1550);
   U3898 : AO4 port map( A => n4207, B => n81, C => n4206, D => n229, Z => 
                           n1551);
   U3899 : AO4 port map( A => n4209, B => n270, C => n4208, D => n272, Z => 
                           n1552);
   U3900 : AO4 port map( A => n4211, B => n72, C => n4210, D => n228, Z => 
                           n1553);
   U3901 : NR4 port map( A => n1555, B => n1556, C => n1557, D => n1558, Z => 
                           n1549);
   U3902 : AO4 port map( A => n4215, B => n71, C => n4214, D => n227, Z => 
                           n1555);
   U3903 : AO4 port map( A => n4217, B => n255, C => n4216, D => n257, Z => 
                           n1556);
   U3904 : AO4 port map( A => n4219, B => n12, C => n4218, D => n23, Z => n1557
                           );
   U3905 : NR4 port map( A => n1559, B => n1560, C => n1561, D => n1562, Z => 
                           n1548);
   U3906 : AO4 port map( A => n4223, B => n69, C => n4222, D => n224, Z => 
                           n1559);
   U3907 : AO4 port map( A => n4225, B => n265, C => n4224, D => n269, Z => 
                           n1560);
   U3908 : AO4 port map( A => n4227, B => n11, C => n4226, D => n217, Z => 
                           n1561);
   U3909 : NR4 port map( A => n1563, B => n1564, C => n1565, D => n1566, Z => 
                           n1547);
   U3910 : AO4 port map( A => n4231, B => n59, C => n4230, D => n209, Z => 
                           n1563);
   U3911 : AO4 port map( A => n4233, B => n251, C => n4232, D => n253, Z => 
                           n1564);
   U3912 : AO4 port map( A => n4235, B => n10, C => n4234, D => n22, Z => n1565
                           );
   U3913 : NR4 port map( A => n1571, B => n1572, C => n1573, D => n1574, Z => 
                           n1570);
   U3914 : AO4 port map( A => n4175, B => n58, C => n4174, D => n200, Z => 
                           n1571);
   U3915 : AO4 port map( A => n4177, B => n260, C => n4176, D => n261, Z => 
                           n1572);
   U3916 : AO4 port map( A => n4179, B => n9, C => n4178, D => n180, Z => n1573
                           );
   U3917 : NR4 port map( A => n1575, B => n1576, C => n1577, D => n1578, Z => 
                           n1569);
   U3918 : AO4 port map( A => n4183, B => n53, C => n4182, D => n170, Z => 
                           n1575);
   U3919 : AO4 port map( A => n4185, B => n249, C => n4184, D => n250, Z => 
                           n1576);
   U3920 : AO4 port map( A => n4187, B => n28, C => n4186, D => n14, Z => n1577
                           );
   U3921 : NR4 port map( A => n1579, B => n1580, C => n1581, D => n1582, Z => 
                           n1568);
   U3922 : AO4 port map( A => n4191, B => n8, C => n4190, D => n163, Z => n1579
                           );
   U3923 : AO4 port map( A => n4193, B => n258, C => n4192, D => n259, Z => 
                           n1580);
   U3924 : AO4 port map( A => n4195, B => n7, C => n4194, D => n150, Z => n1581
                           );
   U3925 : NR4 port map( A => n1583, B => n1584, C => n1585, D => n1586, Z => 
                           n1567);
   U3926 : AO4 port map( A => n4199, B => n48, C => n4198, D => n122, Z => 
                           n1583);
   U3927 : AO4 port map( A => n4201, B => n246, C => n4200, D => n248, Z => 
                           n1584);
   U3928 : AO4 port map( A => n4203, B => n6, C => n4202, D => n109, Z => n1585
                           );
   U3929 : NR4 port map( A => n1595, B => n1596, C => n1597, D => n1598, Z => 
                           n1594);
   U3930 : AO4 port map( A => n4271, B => n81, C => n4270, D => n229, Z => 
                           n1595);
   U3931 : AO4 port map( A => n4273, B => n270, C => n4272, D => n272, Z => 
                           n1596);
   U3932 : AO4 port map( A => n4275, B => n72, C => n4274, D => n228, Z => 
                           n1597);
   U3933 : NR4 port map( A => n1599, B => n1600, C => n1601, D => n1602, Z => 
                           n1593);
   U3934 : AO4 port map( A => n4279, B => n71, C => n4278, D => n227, Z => 
                           n1599);
   U3935 : AO4 port map( A => n4281, B => n255, C => n4280, D => n257, Z => 
                           n1600);
   U3936 : AO4 port map( A => n4283, B => n12, C => n4282, D => n23, Z => n1601
                           );
   U3937 : NR4 port map( A => n1603, B => n1604, C => n1605, D => n1606, Z => 
                           n1592);
   U3938 : AO4 port map( A => n4287, B => n69, C => n4286, D => n224, Z => 
                           n1603);
   U3939 : AO4 port map( A => n4289, B => n265, C => n4288, D => n269, Z => 
                           n1604);
   U3940 : AO4 port map( A => n4291, B => n11, C => n4290, D => n217, Z => 
                           n1605);
   U3941 : NR4 port map( A => n1607, B => n1608, C => n1609, D => n1610, Z => 
                           n1591);
   U3942 : AO4 port map( A => n4295, B => n59, C => n4294, D => n209, Z => 
                           n1607);
   U3943 : AO4 port map( A => n4297, B => n251, C => n4296, D => n253, Z => 
                           n1608);
   U3944 : AO4 port map( A => n4299, B => n10, C => n4298, D => n22, Z => n1609
                           );
   U3945 : NR4 port map( A => n1615, B => n1616, C => n1617, D => n1618, Z => 
                           n1614);
   U3946 : AO4 port map( A => n4239, B => n58, C => n4238, D => n200, Z => 
                           n1615);
   U3947 : AO4 port map( A => n4241, B => n260, C => n4240, D => n261, Z => 
                           n1616);
   U3948 : AO4 port map( A => n4243, B => n9, C => n4242, D => n180, Z => n1617
                           );
   U3949 : NR4 port map( A => n1619, B => n1620, C => n1621, D => n1622, Z => 
                           n1613);
   U3950 : AO4 port map( A => n4247, B => n53, C => n4246, D => n170, Z => 
                           n1619);
   U3951 : AO4 port map( A => n4249, B => n249, C => n4248, D => n250, Z => 
                           n1620);
   U3952 : AO4 port map( A => n4251, B => n28, C => n4250, D => n14, Z => n1621
                           );
   U3953 : NR4 port map( A => n1623, B => n1624, C => n1625, D => n1626, Z => 
                           n1612);
   U3954 : AO4 port map( A => n4255, B => n8, C => n4254, D => n163, Z => n1623
                           );
   U3955 : AO4 port map( A => n4257, B => n258, C => n4256, D => n259, Z => 
                           n1624);
   U3956 : AO4 port map( A => n4259, B => n7, C => n4258, D => n150, Z => n1625
                           );
   U3957 : NR4 port map( A => n1627, B => n1628, C => n1629, D => n1630, Z => 
                           n1611);
   U3958 : AO4 port map( A => n4263, B => n48, C => n4262, D => n122, Z => 
                           n1627);
   U3959 : AO4 port map( A => n4265, B => n246, C => n4264, D => n248, Z => 
                           n1628);
   U3960 : AO4 port map( A => n4267, B => n6, C => n4266, D => n109, Z => n1629
                           );
   U3961 : NR4 port map( A => n1639, B => n1640, C => n1641, D => n1642, Z => 
                           n1638);
   U3962 : AO4 port map( A => n4335, B => n81, C => n4334, D => n229, Z => 
                           n1639);
   U3963 : AO4 port map( A => n4337, B => n270, C => n4336, D => n272, Z => 
                           n1640);
   U3964 : AO4 port map( A => n4339, B => n72, C => n4338, D => n228, Z => 
                           n1641);
   U3965 : NR4 port map( A => n1643, B => n1644, C => n1645, D => n1646, Z => 
                           n1637);
   U3966 : AO4 port map( A => n4343, B => n71, C => n4342, D => n227, Z => 
                           n1643);
   U3967 : AO4 port map( A => n4345, B => n255, C => n4344, D => n257, Z => 
                           n1644);
   U3968 : AO4 port map( A => n4347, B => n12, C => n4346, D => n23, Z => n1645
                           );
   U3969 : NR4 port map( A => n1647, B => n1648, C => n1649, D => n1650, Z => 
                           n1636);
   U3970 : AO4 port map( A => n4351, B => n69, C => n4350, D => n224, Z => 
                           n1647);
   U3971 : AO4 port map( A => n4353, B => n265, C => n4352, D => n269, Z => 
                           n1648);
   U3972 : AO4 port map( A => n4355, B => n11, C => n4354, D => n217, Z => 
                           n1649);
   U3973 : NR4 port map( A => n1651, B => n1652, C => n1653, D => n1654, Z => 
                           n1635);
   U3974 : AO4 port map( A => n4359, B => n59, C => n4358, D => n209, Z => 
                           n1651);
   U3975 : AO4 port map( A => n4361, B => n251, C => n4360, D => n253, Z => 
                           n1652);
   U3976 : AO4 port map( A => n4363, B => n10, C => n4362, D => n22, Z => n1653
                           );
   U3977 : NR4 port map( A => n1659, B => n1660, C => n1661, D => n1662, Z => 
                           n1658);
   U3978 : AO4 port map( A => n4303, B => n58, C => n4302, D => n200, Z => 
                           n1659);
   U3979 : AO4 port map( A => n4305, B => n260, C => n4304, D => n261, Z => 
                           n1660);
   U3980 : AO4 port map( A => n4307, B => n9, C => n4306, D => n180, Z => n1661
                           );
   U3981 : NR4 port map( A => n1663, B => n1664, C => n1665, D => n1666, Z => 
                           n1657);
   U3982 : AO4 port map( A => n4311, B => n53, C => n4310, D => n170, Z => 
                           n1663);
   U3983 : AO4 port map( A => n4313, B => n249, C => n4312, D => n250, Z => 
                           n1664);
   U3984 : AO4 port map( A => n4315, B => n28, C => n4314, D => n14, Z => n1665
                           );
   U3985 : NR4 port map( A => n1667, B => n1668, C => n1669, D => n1670, Z => 
                           n1656);
   U3986 : AO4 port map( A => n4319, B => n8, C => n4318, D => n163, Z => n1667
                           );
   U3987 : AO4 port map( A => n4321, B => n258, C => n4320, D => n259, Z => 
                           n1668);
   U3988 : AO4 port map( A => n4323, B => n7, C => n4322, D => n150, Z => n1669
                           );
   U3989 : NR4 port map( A => n1671, B => n1672, C => n1673, D => n1674, Z => 
                           n1655);
   U3990 : AO4 port map( A => n4327, B => n48, C => n4326, D => n122, Z => 
                           n1671);
   U3991 : AO4 port map( A => n4329, B => n246, C => n4328, D => n248, Z => 
                           n1672);
   U3992 : AO4 port map( A => n4331, B => n6, C => n4330, D => n109, Z => n1673
                           );
   U3993 : NR4 port map( A => n1683, B => n1684, C => n1685, D => n1686, Z => 
                           n1682);
   U3994 : AO4 port map( A => n4399, B => n81, C => n4398, D => n229, Z => 
                           n1683);
   U3995 : AO4 port map( A => n4401, B => n270, C => n4400, D => n272, Z => 
                           n1684);
   U3996 : AO4 port map( A => n4403, B => n72, C => n4402, D => n228, Z => 
                           n1685);
   U3997 : NR4 port map( A => n1687, B => n1688, C => n1689, D => n1690, Z => 
                           n1681);
   U3998 : AO4 port map( A => n4407, B => n71, C => n4406, D => n227, Z => 
                           n1687);
   U3999 : AO4 port map( A => n4409, B => n255, C => n4408, D => n257, Z => 
                           n1688);
   U4000 : AO4 port map( A => n4411, B => n12, C => n4410, D => n23, Z => n1689
                           );
   U4001 : NR4 port map( A => n1691, B => n1692, C => n1693, D => n1694, Z => 
                           n1680);
   U4002 : AO4 port map( A => n4415, B => n69, C => n4414, D => n224, Z => 
                           n1691);
   U4003 : AO4 port map( A => n4417, B => n265, C => n4416, D => n269, Z => 
                           n1692);
   U4004 : AO4 port map( A => n4419, B => n11, C => n4418, D => n217, Z => 
                           n1693);
   U4005 : NR4 port map( A => n1695, B => n1696, C => n1697, D => n1698, Z => 
                           n1679);
   U4006 : AO4 port map( A => n4423, B => n59, C => n4422, D => n209, Z => 
                           n1695);
   U4007 : AO4 port map( A => n4425, B => n251, C => n4424, D => n253, Z => 
                           n1696);
   U4008 : AO4 port map( A => n4427, B => n10, C => n4426, D => n22, Z => n1697
                           );
   U4009 : NR4 port map( A => n1703, B => n1704, C => n1705, D => n1706, Z => 
                           n1702);
   U4010 : AO4 port map( A => n4367, B => n58, C => n4366, D => n200, Z => 
                           n1703);
   U4011 : AO4 port map( A => n4369, B => n260, C => n4368, D => n261, Z => 
                           n1704);
   U4012 : AO4 port map( A => n4371, B => n9, C => n4370, D => n180, Z => n1705
                           );
   U4013 : NR4 port map( A => n1707, B => n1708, C => n1709, D => n1710, Z => 
                           n1701);
   U4014 : AO4 port map( A => n4375, B => n53, C => n4374, D => n170, Z => 
                           n1707);
   U4015 : AO4 port map( A => n4377, B => n249, C => n4376, D => n250, Z => 
                           n1708);
   U4016 : AO4 port map( A => n4379, B => n28, C => n4378, D => n14, Z => n1709
                           );
   U4017 : NR4 port map( A => n1711, B => n1712, C => n1713, D => n1714, Z => 
                           n1700);
   U4018 : AO4 port map( A => n4383, B => n8, C => n4382, D => n163, Z => n1711
                           );
   U4019 : AO4 port map( A => n4385, B => n258, C => n4384, D => n259, Z => 
                           n1712);
   U4020 : AO4 port map( A => n4387, B => n7, C => n4386, D => n150, Z => n1713
                           );
   U4021 : NR4 port map( A => n1715, B => n1716, C => n1717, D => n1718, Z => 
                           n1699);
   U4022 : AO4 port map( A => n4391, B => n48, C => n4390, D => n122, Z => 
                           n1715);
   U4023 : AO4 port map( A => n4393, B => n246, C => n4392, D => n248, Z => 
                           n1716);
   U4024 : AO4 port map( A => n4395, B => n6, C => n4394, D => n109, Z => n1717
                           );
   U4025 : NR4 port map( A => n1727, B => n1728, C => n1729, D => n1730, Z => 
                           n1726);
   U4026 : AO4 port map( A => n4463, B => n81, C => n4462, D => n229, Z => 
                           n1727);
   U4027 : AO4 port map( A => n4465, B => n270, C => n4464, D => n272, Z => 
                           n1728);
   U4028 : AO4 port map( A => n4467, B => n72, C => n4466, D => n228, Z => 
                           n1729);
   U4029 : NR4 port map( A => n1731, B => n1732, C => n1733, D => n1734, Z => 
                           n1725);
   U4030 : AO4 port map( A => n4471, B => n71, C => n4470, D => n227, Z => 
                           n1731);
   U4031 : AO4 port map( A => n4473, B => n255, C => n4472, D => n257, Z => 
                           n1732);
   U4032 : AO4 port map( A => n4475, B => n12, C => n4474, D => n23, Z => n1733
                           );
   U4033 : NR4 port map( A => n1735, B => n1736, C => n1737, D => n1738, Z => 
                           n1724);
   U4034 : AO4 port map( A => n4479, B => n69, C => n4478, D => n224, Z => 
                           n1735);
   U4035 : AO4 port map( A => n4481, B => n265, C => n4480, D => n269, Z => 
                           n1736);
   U4036 : AO4 port map( A => n4483, B => n11, C => n4482, D => n217, Z => 
                           n1737);
   U4037 : NR4 port map( A => n1739, B => n1740, C => n1741, D => n1742, Z => 
                           n1723);
   U4038 : AO4 port map( A => n4487, B => n59, C => n4486, D => n209, Z => 
                           n1739);
   U4039 : AO4 port map( A => n4489, B => n251, C => n4488, D => n253, Z => 
                           n1740);
   U4040 : AO4 port map( A => n4491, B => n10, C => n4490, D => n22, Z => n1741
                           );
   U4041 : NR4 port map( A => n1747, B => n1748_port, C => n1749_port, D => 
                           n1750_port, Z => n1746);
   U4042 : AO4 port map( A => n4431, B => n58, C => n4430, D => n200, Z => 
                           n1747);
   U4043 : AO4 port map( A => n4433, B => n260, C => n4432, D => n261, Z => 
                           n1748_port);
   U4044 : AO4 port map( A => n4435, B => n9, C => n4434, D => n180, Z => 
                           n1749_port);
   U4045 : NR4 port map( A => n1751_port, B => n1752_port, C => n1753_port, D 
                           => n1754_port, Z => n1745);
   U4046 : AO4 port map( A => n4439, B => n53, C => n4438, D => n170, Z => 
                           n1751_port);
   U4047 : AO4 port map( A => n4441, B => n249, C => n4440, D => n250, Z => 
                           n1752_port);
   U4048 : AO4 port map( A => n4443, B => n28, C => n4442, D => n14, Z => 
                           n1753_port);
   U4049 : NR4 port map( A => n1755, B => n1756, C => n1757, D => n1758, Z => 
                           n1744);
   U4050 : AO4 port map( A => n4447, B => n8, C => n4446, D => n163, Z => n1755
                           );
   U4051 : AO4 port map( A => n4449, B => n258, C => n4448, D => n259, Z => 
                           n1756);
   U4052 : AO4 port map( A => n4451, B => n7, C => n4450, D => n150, Z => n1757
                           );
   U4053 : NR4 port map( A => n1759, B => n1760, C => n1761, D => n1762, Z => 
                           n1743);
   U4054 : AO4 port map( A => n4455, B => n48, C => n4454, D => n122, Z => 
                           n1759);
   U4055 : AO4 port map( A => n4457, B => n246, C => n4456, D => n248, Z => 
                           n1760);
   U4056 : AO4 port map( A => n4459, B => n6, C => n4458, D => n109, Z => n1761
                           );
   U4057 : NR4 port map( A => n1771, B => n1772, C => n1773, D => n1774, Z => 
                           n1770);
   U4058 : AO4 port map( A => n4527, B => n81, C => n4526, D => n229, Z => 
                           n1771);
   U4059 : AO4 port map( A => n4529, B => n270, C => n4528, D => n272, Z => 
                           n1772);
   U4060 : AO4 port map( A => n4531, B => n72, C => n4530, D => n228, Z => 
                           n1773);
   U4061 : NR4 port map( A => n1784, B => n1785, C => n1786, D => n1787, Z => 
                           n1769);
   U4062 : AO4 port map( A => n4535, B => n71, C => n4534, D => n227, Z => 
                           n1784);
   U4063 : AO4 port map( A => n4537, B => n255, C => n4536, D => n257, Z => 
                           n1785);
   U4064 : AO4 port map( A => n4539, B => n12, C => n4538, D => n23, Z => n1786
                           );
   U4065 : NR4 port map( A => n1794, B => n1795, C => n1796, D => n1797, Z => 
                           n1768);
   U4066 : AO4 port map( A => n4543, B => n69, C => n4542, D => n224, Z => 
                           n1794);
   U4067 : AO4 port map( A => n4545, B => n265, C => n4544, D => n269, Z => 
                           n1795);
   U4068 : AO4 port map( A => n4547, B => n11, C => n4546, D => n217, Z => 
                           n1796);
   U4069 : NR4 port map( A => n1801, B => n1802, C => n1803, D => n1804, Z => 
                           n1767);
   U4070 : AO4 port map( A => n4551, B => n59, C => n4550, D => n209, Z => 
                           n1801);
   U4071 : AO4 port map( A => n4553, B => n251, C => n4552, D => n253, Z => 
                           n1802);
   U4072 : AO4 port map( A => n4555, B => n10, C => n4554, D => n22, Z => n1803
                           );
   U4073 : NR4 port map( A => n1813, B => n1814, C => n1815, D => n1816, Z => 
                           n1812);
   U4074 : AO4 port map( A => n4495, B => n58, C => n4494, D => n200, Z => 
                           n1813);
   U4075 : AO4 port map( A => n4497, B => n260, C => n4496, D => n261, Z => 
                           n1814);
   U4076 : AO4 port map( A => n4499, B => n9, C => n4498, D => n180, Z => n1815
                           );
   U4077 : NR4 port map( A => n1820, B => n1821, C => n1822, D => n1823, Z => 
                           n1811);
   U4078 : AO4 port map( A => n4503, B => n53, C => n4502, D => n170, Z => 
                           n1820);
   U4079 : AO4 port map( A => n4505, B => n249, C => n4504, D => n250, Z => 
                           n1821);
   U4080 : AO4 port map( A => n4507, B => n28, C => n4506, D => n14, Z => n1822
                           );
   U4081 : NR4 port map( A => n1826, B => n1827, C => n1828, D => n1829, Z => 
                           n1810);
   U4082 : AO4 port map( A => n4511, B => n8, C => n4510, D => n163, Z => n1826
                           );
   U4083 : AO4 port map( A => n4513, B => n258, C => n4512, D => n259, Z => 
                           n1827);
   U4084 : AO4 port map( A => n4515, B => n7, C => n4514, D => n150, Z => n1828
                           );
   U4085 : NR4 port map( A => n1837, B => n1838, C => n1839, D => n1840, Z => 
                           n1809);
   U4086 : AO4 port map( A => n4519, B => n48, C => n4518, D => n122, Z => 
                           n1837);
   U4087 : AO4 port map( A => n4521, B => n246, C => n4520, D => n248, Z => 
                           n1838);
   U4088 : AO4 port map( A => n4523, B => n6, C => n4522, D => n109, Z => n1839
                           );
   U4089 : EON1 port map( A => KEY_NUMB_I(1), B => n6807, C => n6807, D => 
                           n6663, Z => n1846);
   U4090 : EON1 port map( A => KEY_NUMB_I(0), B => n6807, C => n6807, D => 
                           n6664, Z => n1845);
   U4091 : EON1 port map( A => KEY_NUMB_I(2), B => n6807, C => n6807, D => 
                           n6662, Z => n1835);
   U4092 : EON1 port map( A => KEY_NUMB_I(3), B => n6807, C => n6807, D => 
                           n6661, Z => n1836);
   U4093 : EON1 port map( A => KEY_NUMB_I(5), B => n6807, C => n6807, D => 
                           n6659, Z => n1808);
   U4094 : EON1 port map( A => KEY_NUMB_I(4), B => n6807, C => n6807, D => 
                           n6660, Z => n1807);
   U4095 : AO6 port map( A => n6791, B => n6677, C => n287, Z => n283);
   U4096 : IVI port map( A => GET_KEY_I, Z => n6807);
   U4097 : AO4 port map( A => n2549, B => n3, C => n2548, D => n5, Z => n346);
   U4098 : AO4 port map( A => n2557, B => n2, C => n2556, D => n4, Z => n358);
   U4099 : AO4 port map( A => n2565, B => n43, C => n2564, D => n33, Z => n370)
                           ;
   U4100 : AO4 port map( A => n2573, B => n1, C => n2572, D => n38, Z => n382);
   U4101 : AO4 port map( A => n2517, B => n241, C => n2516, D => n245, Z => 
                           n398);
   U4102 : AO4 port map( A => n2525, B => n237, C => n2524, D => n238, Z => 
                           n410);
   U4103 : AO4 port map( A => n2533, B => n235, C => n2532, D => n236, Z => 
                           n422);
   U4104 : AO4 port map( A => n2541, B => n232, C => n2540, D => n234, Z => 
                           n434);
   U4105 : AO4 port map( A => n2613, B => n3, C => n2612, D => n5, Z => n454);
   U4106 : AO4 port map( A => n2621, B => n2, C => n2620, D => n4, Z => n458);
   U4107 : AO4 port map( A => n2629, B => n43, C => n2628, D => n33, Z => n462)
                           ;
   U4108 : AO4 port map( A => n2637, B => n1, C => n2636, D => n38, Z => n466);
   U4109 : AO4 port map( A => n2581, B => n241, C => n2580, D => n245, Z => 
                           n474);
   U4110 : AO4 port map( A => n2589, B => n237, C => n2588, D => n238, Z => 
                           n478);
   U4111 : AO4 port map( A => n2597, B => n235, C => n2596, D => n236, Z => 
                           n482);
   U4112 : AO4 port map( A => n2605, B => n232, C => n2604, D => n234, Z => 
                           n486);
   U4113 : AO4 port map( A => n2677, B => n3, C => n2676, D => n5, Z => n498);
   U4114 : AO4 port map( A => n2685, B => n2, C => n2684, D => n4, Z => n502);
   U4115 : AO4 port map( A => n2693, B => n43, C => n2692, D => n33, Z => n506)
                           ;
   U4116 : AO4 port map( A => n2701, B => n1, C => n2700, D => n38, Z => n510);
   U4117 : AO4 port map( A => n2645, B => n241, C => n2644, D => n245, Z => 
                           n518);
   U4118 : AO4 port map( A => n2653, B => n237, C => n2652, D => n238, Z => 
                           n522);
   U4119 : AO4 port map( A => n2661, B => n235, C => n2660, D => n236, Z => 
                           n526);
   U4120 : AO4 port map( A => n2669, B => n232, C => n2668, D => n234, Z => 
                           n530);
   U4121 : AO4 port map( A => n2741, B => n3, C => n2740, D => n5, Z => n542);
   U4122 : AO4 port map( A => n2749, B => n2, C => n2748, D => n4, Z => n546);
   U4123 : AO4 port map( A => n2757, B => n43, C => n2756, D => n33, Z => n550)
                           ;
   U4124 : AO4 port map( A => n2765, B => n1, C => n2764, D => n38, Z => n554);
   U4125 : AO4 port map( A => n2709, B => n241, C => n2708, D => n245, Z => 
                           n562);
   U4126 : AO4 port map( A => n2717, B => n237, C => n2716, D => n238, Z => 
                           n566);
   U4127 : AO4 port map( A => n2725, B => n235, C => n2724, D => n236, Z => 
                           n570);
   U4128 : AO4 port map( A => n2733, B => n232, C => n2732, D => n234, Z => 
                           n574);
   U4129 : AO4 port map( A => n2805, B => n3, C => n2804, D => n5, Z => n586);
   U4130 : AO4 port map( A => n2813, B => n2, C => n2812, D => n4, Z => n590);
   U4131 : AO4 port map( A => n2821, B => n43, C => n2820, D => n33, Z => n594)
                           ;
   U4132 : AO4 port map( A => n2829, B => n1, C => n2828, D => n38, Z => n598);
   U4133 : AO4 port map( A => n2773, B => n241, C => n2772, D => n245, Z => 
                           n606);
   U4134 : AO4 port map( A => n2781, B => n237, C => n2780, D => n238, Z => 
                           n610);
   U4135 : AO4 port map( A => n2789, B => n235, C => n2788, D => n236, Z => 
                           n614);
   U4136 : AO4 port map( A => n2797, B => n232, C => n2796, D => n234, Z => 
                           n618);
   U4137 : AO4 port map( A => n2869, B => n3, C => n2868, D => n5, Z => n630);
   U4138 : AO4 port map( A => n2877, B => n2, C => n2876, D => n4, Z => n634);
   U4139 : AO4 port map( A => n2885, B => n43, C => n2884, D => n33, Z => n638)
                           ;
   U4140 : AO4 port map( A => n2893, B => n1, C => n2892, D => n38, Z => n642);
   U4141 : AO4 port map( A => n2837, B => n241, C => n2836, D => n245, Z => 
                           n650);
   U4142 : AO4 port map( A => n2845, B => n237, C => n2844, D => n238, Z => 
                           n654);
   U4143 : AO4 port map( A => n2853, B => n235, C => n2852, D => n236, Z => 
                           n658);
   U4144 : AO4 port map( A => n2861, B => n232, C => n2860, D => n234, Z => 
                           n662);
   U4145 : AO4 port map( A => n2933, B => n3, C => n2932, D => n5, Z => n674);
   U4146 : AO4 port map( A => n2941, B => n2, C => n2940, D => n4, Z => n678);
   U4147 : AO4 port map( A => n2949, B => n43, C => n2948, D => n33, Z => n682)
                           ;
   U4148 : AO4 port map( A => n2957, B => n1, C => n2956, D => n38, Z => n686);
   U4149 : AO4 port map( A => n2901, B => n241, C => n2900, D => n245, Z => 
                           n694);
   U4150 : AO4 port map( A => n2909, B => n237, C => n2908, D => n238, Z => 
                           n698);
   U4151 : AO4 port map( A => n2917, B => n235, C => n2916, D => n236, Z => 
                           n702);
   U4152 : AO4 port map( A => n2925, B => n232, C => n2924, D => n234, Z => 
                           n706);
   U4153 : AO4 port map( A => n2997, B => n3, C => n2996, D => n5, Z => n718);
   U4154 : AO4 port map( A => n3005, B => n2, C => n3004, D => n4, Z => n722);
   U4155 : AO4 port map( A => n3013, B => n43, C => n3012, D => n33, Z => n726)
                           ;
   U4156 : AO4 port map( A => n3021, B => n1, C => n3020, D => n38, Z => n730);
   U4157 : AO4 port map( A => n2965, B => n241, C => n2964, D => n245, Z => 
                           n738);
   U4158 : AO4 port map( A => n2973, B => n237, C => n2972, D => n238, Z => 
                           n742);
   U4159 : AO4 port map( A => n2981, B => n235, C => n2980, D => n236, Z => 
                           n746);
   U4160 : AO4 port map( A => n2989, B => n232, C => n2988, D => n234, Z => 
                           n750);
   U4161 : AO4 port map( A => n3061, B => n3, C => n3060, D => n5, Z => n762);
   U4162 : AO4 port map( A => n3069, B => n2, C => n3068, D => n4, Z => n766);
   U4163 : AO4 port map( A => n3077, B => n43, C => n3076, D => n33, Z => n770)
                           ;
   U4164 : AO4 port map( A => n3085, B => n1, C => n3084, D => n38, Z => n774);
   U4165 : AO4 port map( A => n3029, B => n241, C => n3028, D => n245, Z => 
                           n782);
   U4166 : AO4 port map( A => n3037, B => n237, C => n3036, D => n238, Z => 
                           n786);
   U4167 : AO4 port map( A => n3045, B => n235, C => n3044, D => n236, Z => 
                           n790);
   U4168 : AO4 port map( A => n3053, B => n232, C => n3052, D => n234, Z => 
                           n794);
   U4169 : AO4 port map( A => n3125, B => n3, C => n3124, D => n5, Z => n806);
   U4170 : AO4 port map( A => n3133, B => n2, C => n3132, D => n4, Z => n810);
   U4171 : AO4 port map( A => n3141, B => n43, C => n3140, D => n33, Z => n814)
                           ;
   U4172 : AO4 port map( A => n3149, B => n1, C => n3148, D => n38, Z => n818);
   U4173 : AO4 port map( A => n3093, B => n241, C => n3092, D => n245, Z => 
                           n826);
   U4174 : AO4 port map( A => n3101, B => n237, C => n3100, D => n238, Z => 
                           n830);
   U4175 : AO4 port map( A => n3109, B => n235, C => n3108, D => n236, Z => 
                           n834);
   U4176 : AO4 port map( A => n3117, B => n232, C => n3116, D => n234, Z => 
                           n838);
   U4177 : AO4 port map( A => n3189, B => n3, C => n3188, D => n5, Z => n850);
   U4178 : AO4 port map( A => n3197, B => n2, C => n3196, D => n4, Z => n854);
   U4179 : AO4 port map( A => n3205, B => n43, C => n3204, D => n33, Z => n858)
                           ;
   U4180 : AO4 port map( A => n3213, B => n1, C => n3212, D => n38, Z => n862);
   U4181 : AO4 port map( A => n3157, B => n241, C => n3156, D => n245, Z => 
                           n870);
   U4182 : AO4 port map( A => n3165, B => n237, C => n3164, D => n238, Z => 
                           n874);
   U4183 : AO4 port map( A => n3173, B => n235, C => n3172, D => n236, Z => 
                           n878);
   U4184 : AO4 port map( A => n3181, B => n232, C => n3180, D => n234, Z => 
                           n882);
   U4185 : AO4 port map( A => n3253, B => n3, C => n3252, D => n5, Z => n894);
   U4186 : AO4 port map( A => n3261, B => n2, C => n3260, D => n4, Z => n898);
   U4187 : AO4 port map( A => n3269, B => n43, C => n3268, D => n33, Z => n902)
                           ;
   U4188 : AO4 port map( A => n3277, B => n1, C => n3276, D => n38, Z => n906);
   U4189 : AO4 port map( A => n3221, B => n241, C => n3220, D => n245, Z => 
                           n914);
   U4190 : AO4 port map( A => n3229, B => n237, C => n3228, D => n238, Z => 
                           n918);
   U4191 : AO4 port map( A => n3237, B => n235, C => n3236, D => n236, Z => 
                           n922);
   U4192 : AO4 port map( A => n3245, B => n232, C => n3244, D => n234, Z => 
                           n926);
   U4193 : AO4 port map( A => n3317, B => n3, C => n3316, D => n5, Z => n938);
   U4194 : AO4 port map( A => n3325, B => n2, C => n3324, D => n4, Z => n942);
   U4195 : AO4 port map( A => n3333, B => n43, C => n3332, D => n33, Z => n946)
                           ;
   U4196 : AO4 port map( A => n3341, B => n1, C => n3340, D => n38, Z => n950);
   U4197 : AO4 port map( A => n3285, B => n241, C => n3284, D => n245, Z => 
                           n958);
   U4198 : AO4 port map( A => n3293, B => n237, C => n3292, D => n238, Z => 
                           n962);
   U4199 : AO4 port map( A => n3301, B => n235, C => n3300, D => n236, Z => 
                           n966);
   U4200 : AO4 port map( A => n3309, B => n232, C => n3308, D => n234, Z => 
                           n970);
   U4201 : AO4 port map( A => n3381, B => n3, C => n3380, D => n5, Z => n982);
   U4202 : AO4 port map( A => n3389, B => n2, C => n3388, D => n4, Z => n986);
   U4203 : AO4 port map( A => n3397, B => n43, C => n3396, D => n33, Z => n990)
                           ;
   U4204 : AO4 port map( A => n3405, B => n1, C => n3404, D => n38, Z => n994);
   U4205 : AO4 port map( A => n3349, B => n241, C => n3348, D => n245, Z => 
                           n1002);
   U4206 : AO4 port map( A => n3357, B => n237, C => n3356, D => n238, Z => 
                           n1006);
   U4207 : AO4 port map( A => n3365, B => n235, C => n3364, D => n236, Z => 
                           n1010);
   U4208 : AO4 port map( A => n3373, B => n232, C => n3372, D => n234, Z => 
                           n1014);
   U4209 : AO4 port map( A => n3445, B => n3, C => n3444, D => n5, Z => n1026);
   U4210 : AO4 port map( A => n3453, B => n2, C => n3452, D => n4, Z => n1030);
   U4211 : AO4 port map( A => n3461, B => n43, C => n3460, D => n33, Z => n1034
                           );
   U4212 : AO4 port map( A => n3469, B => n1, C => n3468, D => n38, Z => n1038)
                           ;
   U4213 : AO4 port map( A => n3413, B => n241, C => n3412, D => n245, Z => 
                           n1046);
   U4214 : AO4 port map( A => n3421, B => n237, C => n3420, D => n238, Z => 
                           n1050);
   U4215 : AO4 port map( A => n3429, B => n235, C => n3428, D => n236, Z => 
                           n1054);
   U4216 : AO4 port map( A => n3437, B => n232, C => n3436, D => n234, Z => 
                           n1058);
   U4217 : AO4 port map( A => n3509, B => n3, C => n3508, D => n5, Z => n1070);
   U4218 : AO4 port map( A => n3517, B => n2, C => n3516, D => n4, Z => n1074);
   U4219 : AO4 port map( A => n3525, B => n43, C => n3524, D => n33, Z => n1078
                           );
   U4220 : AO4 port map( A => n3533, B => n1, C => n3532, D => n38, Z => n1082)
                           ;
   U4221 : AO4 port map( A => n3477, B => n241, C => n3476, D => n245, Z => 
                           n1090);
   U4222 : AO4 port map( A => n3485, B => n237, C => n3484, D => n238, Z => 
                           n1094);
   U4223 : AO4 port map( A => n3493, B => n235, C => n3492, D => n236, Z => 
                           n1098);
   U4224 : AO4 port map( A => n3501, B => n232, C => n3500, D => n234, Z => 
                           n1102);
   U4225 : AO4 port map( A => n3573, B => n3, C => n3572, D => n5, Z => n1114);
   U4226 : AO4 port map( A => n3581, B => n2, C => n3580, D => n4, Z => n1118);
   U4227 : AO4 port map( A => n3589, B => n43, C => n3588, D => n33, Z => n1122
                           );
   U4228 : AO4 port map( A => n3597, B => n1, C => n3596, D => n38, Z => n1126)
                           ;
   U4229 : AO4 port map( A => n3541, B => n241, C => n3540, D => n245, Z => 
                           n1134);
   U4230 : AO4 port map( A => n3549, B => n237, C => n3548, D => n238, Z => 
                           n1138);
   U4231 : AO4 port map( A => n3557, B => n235, C => n3556, D => n236, Z => 
                           n1142);
   U4232 : AO4 port map( A => n3565, B => n232, C => n3564, D => n234, Z => 
                           n1146);
   U4233 : AO4 port map( A => n3637, B => n3, C => n3636, D => n5, Z => n1158);
   U4234 : AO4 port map( A => n3645, B => n2, C => n3644, D => n4, Z => n1162);
   U4235 : AO4 port map( A => n3653, B => n43, C => n3652, D => n33, Z => n1166
                           );
   U4236 : AO4 port map( A => n3661, B => n1, C => n3660, D => n38, Z => n1170)
                           ;
   U4237 : AO4 port map( A => n3605, B => n241, C => n3604, D => n245, Z => 
                           n1178);
   U4238 : AO4 port map( A => n3613, B => n237, C => n3612, D => n238, Z => 
                           n1182);
   U4239 : AO4 port map( A => n3621, B => n235, C => n3620, D => n236, Z => 
                           n1186);
   U4240 : AO4 port map( A => n3629, B => n232, C => n3628, D => n234, Z => 
                           n1190);
   U4241 : AO4 port map( A => n3701, B => n3, C => n3700, D => n5, Z => n1202);
   U4242 : AO4 port map( A => n3709, B => n2, C => n3708, D => n4, Z => n1206);
   U4243 : AO4 port map( A => n3717, B => n43, C => n3716, D => n33, Z => n1210
                           );
   U4244 : AO4 port map( A => n3725, B => n1, C => n3724, D => n38, Z => n1214)
                           ;
   U4245 : AO4 port map( A => n3669, B => n241, C => n3668, D => n245, Z => 
                           n1222);
   U4246 : AO4 port map( A => n3677, B => n237, C => n3676, D => n238, Z => 
                           n1226);
   U4247 : AO4 port map( A => n3685, B => n235, C => n3684, D => n236, Z => 
                           n1230);
   U4248 : AO4 port map( A => n3693, B => n232, C => n3692, D => n234, Z => 
                           n1234);
   U4249 : AO4 port map( A => n3765, B => n3, C => n3764, D => n5, Z => n1246);
   U4250 : AO4 port map( A => n3773, B => n2, C => n3772, D => n4, Z => n1250);
   U4251 : AO4 port map( A => n3781, B => n43, C => n3780, D => n33, Z => n1254
                           );
   U4252 : AO4 port map( A => n3789, B => n1, C => n3788, D => n38, Z => n1258)
                           ;
   U4253 : AO4 port map( A => n3733, B => n241, C => n3732, D => n245, Z => 
                           n1266);
   U4254 : AO4 port map( A => n3741, B => n237, C => n3740, D => n238, Z => 
                           n1270);
   U4255 : AO4 port map( A => n3749, B => n235, C => n3748, D => n236, Z => 
                           n1274);
   U4256 : AO4 port map( A => n3757, B => n232, C => n3756, D => n234, Z => 
                           n1278);
   U4257 : AO4 port map( A => n3829, B => n3, C => n3828, D => n5, Z => n1290);
   U4258 : AO4 port map( A => n3837, B => n2, C => n3836, D => n4, Z => n1294);
   U4259 : AO4 port map( A => n3845, B => n43, C => n3844, D => n33, Z => n1298
                           );
   U4260 : AO4 port map( A => n3853, B => n1, C => n3852, D => n38, Z => n1302)
                           ;
   U4261 : AO4 port map( A => n3797, B => n241, C => n3796, D => n245, Z => 
                           n1310);
   U4262 : AO4 port map( A => n3805, B => n237, C => n3804, D => n238, Z => 
                           n1314);
   U4263 : AO4 port map( A => n3813, B => n235, C => n3812, D => n236, Z => 
                           n1318);
   U4264 : AO4 port map( A => n3821, B => n232, C => n3820, D => n234, Z => 
                           n1322);
   U4265 : AO4 port map( A => n3893, B => n3, C => n3892, D => n5, Z => n1334);
   U4266 : AO4 port map( A => n3901, B => n2, C => n3900, D => n4, Z => n1338);
   U4267 : AO4 port map( A => n3909, B => n43, C => n3908, D => n33, Z => n1342
                           );
   U4268 : AO4 port map( A => n3917, B => n1, C => n3916, D => n38, Z => n1346)
                           ;
   U4269 : AO4 port map( A => n3861, B => n241, C => n3860, D => n245, Z => 
                           n1354);
   U4270 : AO4 port map( A => n3869, B => n237, C => n3868, D => n238, Z => 
                           n1358);
   U4271 : AO4 port map( A => n3877, B => n235, C => n3876, D => n236, Z => 
                           n1362);
   U4272 : AO4 port map( A => n3885, B => n232, C => n3884, D => n234, Z => 
                           n1366);
   U4273 : AO4 port map( A => n3957, B => n3, C => n3956, D => n5, Z => n1378);
   U4274 : AO4 port map( A => n3965, B => n2, C => n3964, D => n4, Z => n1382);
   U4275 : AO4 port map( A => n3973, B => n43, C => n3972, D => n33, Z => n1386
                           );
   U4276 : AO4 port map( A => n3981, B => n1, C => n3980, D => n38, Z => n1390)
                           ;
   U4277 : AO4 port map( A => n3925, B => n241, C => n3924, D => n245, Z => 
                           n1398);
   U4278 : AO4 port map( A => n3933, B => n237, C => n3932, D => n238, Z => 
                           n1402);
   U4279 : AO4 port map( A => n3941, B => n235, C => n3940, D => n236, Z => 
                           n1406);
   U4280 : AO4 port map( A => n3949, B => n232, C => n3948, D => n234, Z => 
                           n1410);
   U4281 : AO4 port map( A => n4021, B => n3, C => n4020, D => n5, Z => n1422);
   U4282 : AO4 port map( A => n4029, B => n2, C => n4028, D => n4, Z => n1426);
   U4283 : AO4 port map( A => n4037, B => n43, C => n4036, D => n33, Z => n1430
                           );
   U4284 : AO4 port map( A => n4045, B => n1, C => n4044, D => n38, Z => n1434)
                           ;
   U4285 : AO4 port map( A => n3989, B => n241, C => n3988, D => n245, Z => 
                           n1442);
   U4286 : AO4 port map( A => n3997, B => n237, C => n3996, D => n238, Z => 
                           n1446);
   U4287 : AO4 port map( A => n4005, B => n235, C => n4004, D => n236, Z => 
                           n1450);
   U4288 : AO4 port map( A => n4013, B => n232, C => n4012, D => n234, Z => 
                           n1454);
   U4289 : AO4 port map( A => n4085, B => n3, C => n4084, D => n5, Z => n1466);
   U4290 : AO4 port map( A => n4093, B => n2, C => n4092, D => n4, Z => n1470);
   U4291 : AO4 port map( A => n4101, B => n43, C => n4100, D => n33, Z => n1474
                           );
   U4292 : AO4 port map( A => n4109, B => n1, C => n4108, D => n38, Z => n1478)
                           ;
   U4293 : AO4 port map( A => n4053, B => n241, C => n4052, D => n245, Z => 
                           n1486);
   U4294 : AO4 port map( A => n4061, B => n237, C => n4060, D => n238, Z => 
                           n1490);
   U4295 : AO4 port map( A => n4069, B => n235, C => n4068, D => n236, Z => 
                           n1494);
   U4296 : AO4 port map( A => n4077, B => n232, C => n4076, D => n234, Z => 
                           n1498);
   U4297 : AO4 port map( A => n4149, B => n3, C => n4148, D => n5, Z => n1510);
   U4298 : AO4 port map( A => n4157, B => n2, C => n4156, D => n4, Z => n1514);
   U4299 : AO4 port map( A => n4165, B => n43, C => n4164, D => n33, Z => n1518
                           );
   U4300 : AO4 port map( A => n4173, B => n1, C => n4172, D => n38, Z => n1522)
                           ;
   U4301 : AO4 port map( A => n4117, B => n241, C => n4116, D => n245, Z => 
                           n1530);
   U4302 : AO4 port map( A => n4125, B => n237, C => n4124, D => n238, Z => 
                           n1534);
   U4303 : AO4 port map( A => n4133, B => n235, C => n4132, D => n236, Z => 
                           n1538);
   U4304 : AO4 port map( A => n4141, B => n232, C => n4140, D => n234, Z => 
                           n1542);
   U4305 : AO4 port map( A => n4213, B => n3, C => n4212, D => n5, Z => n1554);
   U4306 : AO4 port map( A => n4221, B => n2, C => n4220, D => n4, Z => n1558);
   U4307 : AO4 port map( A => n4229, B => n43, C => n4228, D => n33, Z => n1562
                           );
   U4308 : AO4 port map( A => n4237, B => n1, C => n4236, D => n38, Z => n1566)
                           ;
   U4309 : AO4 port map( A => n4181, B => n241, C => n4180, D => n245, Z => 
                           n1574);
   U4310 : AO4 port map( A => n4189, B => n237, C => n4188, D => n238, Z => 
                           n1578);
   U4311 : AO4 port map( A => n4197, B => n235, C => n4196, D => n236, Z => 
                           n1582);
   U4312 : AO4 port map( A => n4205, B => n232, C => n4204, D => n234, Z => 
                           n1586);
   U4313 : AO4 port map( A => n4277, B => n3, C => n4276, D => n5, Z => n1598);
   U4314 : AO4 port map( A => n4285, B => n2, C => n4284, D => n4, Z => n1602);
   U4315 : AO4 port map( A => n4293, B => n43, C => n4292, D => n33, Z => n1606
                           );
   U4316 : AO4 port map( A => n4301, B => n1, C => n4300, D => n38, Z => n1610)
                           ;
   U4317 : AO4 port map( A => n4245, B => n241, C => n4244, D => n245, Z => 
                           n1618);
   U4318 : AO4 port map( A => n4253, B => n237, C => n4252, D => n238, Z => 
                           n1622);
   U4319 : AO4 port map( A => n4261, B => n235, C => n4260, D => n236, Z => 
                           n1626);
   U4320 : AO4 port map( A => n4269, B => n232, C => n4268, D => n234, Z => 
                           n1630);
   U4321 : AO4 port map( A => n4341, B => n3, C => n4340, D => n5, Z => n1642);
   U4322 : AO4 port map( A => n4349, B => n2, C => n4348, D => n4, Z => n1646);
   U4323 : AO4 port map( A => n4357, B => n43, C => n4356, D => n33, Z => n1650
                           );
   U4324 : AO4 port map( A => n4365, B => n1, C => n4364, D => n38, Z => n1654)
                           ;
   U4325 : AO4 port map( A => n4309, B => n241, C => n4308, D => n245, Z => 
                           n1662);
   U4326 : AO4 port map( A => n4317, B => n237, C => n4316, D => n238, Z => 
                           n1666);
   U4327 : AO4 port map( A => n4325, B => n235, C => n4324, D => n236, Z => 
                           n1670);
   U4328 : AO4 port map( A => n4333, B => n232, C => n4332, D => n234, Z => 
                           n1674);
   U4329 : AO4 port map( A => n4405, B => n3, C => n4404, D => n5, Z => n1686);
   U4330 : AO4 port map( A => n4413, B => n2, C => n4412, D => n4, Z => n1690);
   U4331 : AO4 port map( A => n4421, B => n43, C => n4420, D => n33, Z => n1694
                           );
   U4332 : AO4 port map( A => n4429, B => n1, C => n4428, D => n38, Z => n1698)
                           ;
   U4333 : AO4 port map( A => n4373, B => n241, C => n4372, D => n245, Z => 
                           n1706);
   U4334 : AO4 port map( A => n4381, B => n237, C => n4380, D => n238, Z => 
                           n1710);
   U4335 : AO4 port map( A => n4389, B => n235, C => n4388, D => n236, Z => 
                           n1714);
   U4336 : AO4 port map( A => n4397, B => n232, C => n4396, D => n234, Z => 
                           n1718);
   U4337 : AO4 port map( A => n4469, B => n3, C => n4468, D => n5, Z => n1730);
   U4338 : AO4 port map( A => n4477, B => n2, C => n4476, D => n4, Z => n1734);
   U4339 : AO4 port map( A => n4485, B => n43, C => n4484, D => n33, Z => n1738
                           );
   U4340 : AO4 port map( A => n4493, B => n1, C => n4492, D => n38, Z => n1742)
                           ;
   U4341 : AO4 port map( A => n4437, B => n241, C => n4436, D => n245, Z => 
                           n1750_port);
   U4342 : AO4 port map( A => n4445, B => n237, C => n4444, D => n238, Z => 
                           n1754_port);
   U4343 : AO4 port map( A => n4453, B => n235, C => n4452, D => n236, Z => 
                           n1758);
   U4344 : AO4 port map( A => n4461, B => n232, C => n4460, D => n234, Z => 
                           n1762);
   U4345 : AO4 port map( A => n4533, B => n3, C => n4532, D => n5, Z => n1774);
   U4346 : AO4 port map( A => n4541, B => n2, C => n4540, D => n4, Z => n1787);
   U4347 : AO4 port map( A => n4549, B => n43, C => n4548, D => n33, Z => n1797
                           );
   U4348 : AO4 port map( A => n4557, B => n1, C => n4556, D => n38, Z => n1804)
                           ;
   U4349 : AO4 port map( A => n4501, B => n241, C => n4500, D => n245, Z => 
                           n1816);
   U4350 : AO4 port map( A => n4509, B => n237, C => n4508, D => n238, Z => 
                           n1823);
   U4351 : AO4 port map( A => n4517, B => n235, C => n4516, D => n236, Z => 
                           n1829);
   U4352 : AO4 port map( A => n4525, B => n232, C => n4524, D => n234, Z => 
                           n1840);
   U4353 : AO4 port map( A => n6659, B => n254, C => n2098, D => n256, Z => 
                           n6717);
   U4354 : AO4 port map( A => n6660, B => n254, C => n2127, D => n256, Z => 
                           n6718);
   U4355 : AO4 port map( A => n6661, B => n254, C => n2134, D => n256, Z => 
                           n6719);
   U4356 : AO4 port map( A => n6662, B => n254, C => n2175, D => n256, Z => 
                           n6720);
   U4357 : EOI port map( A => n6663, B => i_INTERN_ADDR_RD05, Z => n2274);
   U4358 : AO4 port map( A => n6664, B => n254, C => i_INTERN_ADDR_RD05, D => 
                           n256, Z => n6722);
   U4359 : AO7 port map( A => n65, B => n187, C => n281, Z => n6726);
   U4360 : EO1 port map( A => n201, B => n282, C => n283, D => n6675, Z => n281
                           );
   U4361 : AO7 port map( A => n6673, B => n2391, C => n6806, Z => n155);
   U4362 : AO4 port map( A => n2304, B => n2205, C => n214, D => n168, Z => 
                           n213);
   U4363 : AO4 port map( A => n2304, B => n2217, C => n206, D => n168, Z => 
                           n205);
   U4364 : AO4 port map( A => n2304, B => n2220, C => n198, D => n168, Z => 
                           n197);
   U4365 : AO4 port map( A => n2304, B => n2244, C => n192, D => n168, Z => 
                           n191);
   U4366 : AO4 port map( A => n2304, B => n2233, C => n185, D => n168, Z => 
                           n184);
   U4367 : AO4 port map( A => n2304, B => n2240, C => n167, D => n168, Z => 
                           n165);
   U4368 : EON1 port map( A => n1844, B => n242, C => N1751, D => n2499, Z => 
                           n6669);
   U4369 : EON1 port map( A => n1883, B => n242, C => N1750, D => n2499, Z => 
                           n6668);
   U4370 : EON1 port map( A => n1877, B => n242, C => N1749, D => n2499, Z => 
                           n6667);
   U4371 : EOI port map( A => v_CALCULATION_CNTR_1_port, B => 
                           v_CALCULATION_CNTR_0_port, Z => N1748);
   U4372 : AO4 port map( A => n6676, B => n283, C => n6788, D => n285, Z => 
                           n6727);
   U4373 : AO4 port map( A => n6674, B => n288, C => n6788, D => n289, Z => 
                           n6729);
   U4374 : AO6 port map( A => n6791, B => n6792, C => n287, Z => n288);
   U4375 : EON1 port map( A => n2255, B => n242, C => n2255, D => n2499, Z => 
                           n6665);
   U4376 : NR3 port map( A => n2480, B => n6655, C => i_SRAM_ADDR_WR01, Z => 
                           n2482);
   U4377 : NR3 port map( A => n2480, B => n6654, C => i_SRAM_ADDR_WR02, Z => 
                           n2483);
   U4378 : NR3 port map( A => i_SRAM_ADDR_WR05, B => n6656, C => 
                           i_SRAM_ADDR_WR04, Z => n2475);
   U4379 : NR3 port map( A => n6658, B => n6656, C => i_SRAM_ADDR_WR04, Z => 
                           n2476);
   U4380 : NR3 port map( A => n6657, B => n6656, C => i_SRAM_ADDR_WR05, Z => 
                           n2477);
   U4381 : NR3 port map( A => n1875, B => n1833, C => n2050, Z => n223);
   U4382 : AO2 port map( A => n6805, B => v_CALCULATION_CNTR_7_port, C => N1754
                           , D => n2499, Z => n2503);
   U4383 : AO2 port map( A => n6805, B => v_CALCULATION_CNTR_6_port, C => N1753
                           , D => n2499, Z => n2502);
   U4384 : AO2 port map( A => n6805, B => v_CALCULATION_CNTR_5_port, C => N1752
                           , D => n2499, Z => n2500);
   U4385 : NR3 port map( A => n6655, B => n6654, C => n2480, Z => n2484);
   U4386 : NR3 port map( A => n6656, B => n6657, C => n6658, Z => n2478);
   U4387 : AO6 port map( A => n263, B => n4563, C => RESET_I, Z => n240);
   U4388 : AO7 port map( A => n2509, B => n242, C => n243, Z => n6716);
   U4389 : AO3 port map( A => n157, B => n244, C => n6806, D => CE_I, Z => n243
                           );
   U4390 : AO4 port map( A => v_CALCULATION_CNTR_2_port, B => n230, C => n6804,
                           D => n247, Z => n244);
   U4391 : AO2 port map( A => n2324, B => KEY_I(0), C => n2041, D => 
                           v_KEY32_IN_0_port, Z => n291);
   U4392 : AO2 port map( A => n2324, B => KEY_I(1), C => n2041, D => 
                           v_KEY32_IN_1_port, Z => n294);
   U4393 : AO2 port map( A => n2324, B => KEY_I(2), C => n2041, D => 
                           v_KEY32_IN_2_port, Z => n295);
   U4394 : AO2 port map( A => n2324, B => KEY_I(3), C => n2041, D => 
                           v_KEY32_IN_3_port, Z => n296);
   U4395 : AO2 port map( A => n2324, B => KEY_I(4), C => n2041, D => 
                           v_KEY32_IN_4_port, Z => n297);
   U4396 : AO2 port map( A => n2324, B => KEY_I(5), C => n2041, D => 
                           v_KEY32_IN_5_port, Z => n298);
   U4397 : AO2 port map( A => n2324, B => KEY_I(6), C => n2041, D => 
                           v_KEY32_IN_6_port, Z => n299);
   U4398 : AO2 port map( A => n2324, B => KEY_I(7), C => n2041, D => 
                           v_KEY32_IN_7_port, Z => n300);
   U4399 : NR3 port map( A => n6676, B => n6677, C => n2050, Z => n201);
   U4400 : NR3 port map( A => n6675, B => n6676, C => n6677, Z => n169);
   U4401 : AO6 port map( A => n2506, B => n2505, C => n6803, Z => n312);
   U4402 : AO2 port map( A => n6677, B => n208, C => n6674, D => n1833, Z => 
                           n207);
   U4403 : AO6 port map( A => n2091, B => n6677, C => n201, Z => n199);
   U4404 : AO7 port map( A => n1833, B => n187, C => n6674, Z => n193);
   U4405 : AO4 port map( A => n2507, B => n268, C => n2481, D => n273, Z => 
                           n6724);
   U4406 : AO4 port map( A => n6673, B => n277, C => n2479, D => n278, Z => 
                           n6725);
   U4407 : AO7 port map( A => n6792, B => n2091, C => CE_I, Z => n280);
   U4408 : AO4 port map( A => n6653, B => n231, C => n2101, D => n233, Z => 
                           n6715);
   U4409 : ND3 port map( A => n1833, B => n6676, C => n6675, Z => n216);
   U4410 : AO2 port map( A => KEY_I(0), B => n2076, C => n2323, D => 
                           v_KEY32_IN_8_port, Z => n302);
   U4411 : AO2 port map( A => KEY_I(1), B => n2076, C => n2323, D => 
                           v_KEY32_IN_9_port, Z => n305);
   U4412 : AO2 port map( A => KEY_I(2), B => n2076, C => n2323, D => 
                           v_KEY32_IN_10_port, Z => n306);
   U4413 : AO2 port map( A => KEY_I(3), B => n2076, C => n2323, D => 
                           v_KEY32_IN_11_port, Z => n307);
   U4414 : AO2 port map( A => KEY_I(4), B => n2076, C => n2323, D => 
                           v_KEY32_IN_12_port, Z => n308);
   U4415 : AO2 port map( A => KEY_I(5), B => n2076, C => n2323, D => 
                           v_KEY32_IN_13_port, Z => n309);
   U4416 : AO2 port map( A => KEY_I(6), B => n2076, C => n2323, D => 
                           v_KEY32_IN_14_port, Z => n310);
   U4417 : AO2 port map( A => KEY_I(7), B => n2076, C => n2323, D => 
                           v_KEY32_IN_15_port, Z => n311);
   U4418 : AO2 port map( A => KEY_I(0), B => n2326, C => n2066, D => 
                           v_KEY32_IN_24_port, Z => n323);
   U4419 : AO2 port map( A => KEY_I(1), B => n2326, C => n2066, D => 
                           v_KEY32_IN_25_port, Z => n326);
   U4420 : AO2 port map( A => KEY_I(2), B => n2326, C => n2066, D => 
                           v_KEY32_IN_26_port, Z => n327);
   U4421 : AO2 port map( A => KEY_I(3), B => n2326, C => n2066, D => 
                           v_KEY32_IN_27_port, Z => n328);
   U4422 : AO2 port map( A => KEY_I(4), B => n2326, C => n2066, D => 
                           v_KEY32_IN_28_port, Z => n329);
   U4423 : AO2 port map( A => KEY_I(5), B => n324, C => n2066, D => 
                           v_KEY32_IN_29_port, Z => n330);
   U4424 : AO2 port map( A => KEY_I(6), B => n324, C => n2066, D => 
                           v_KEY32_IN_30_port, Z => n331);
   U4425 : AO2 port map( A => KEY_I(7), B => n324, C => n2066, D => 
                           v_KEY32_IN_31_port, Z => n332);
   U4426 : AO6 port map( A => CE_I, B => n279, C => RESET_I, Z => n274);
   U4427 : AO6 port map( A => n187, B => n6674, C => n6677, Z => n186);
   U4428 : AO4 port map( A => n6654, B => n231, C => n2146, D => n233, Z => 
                           n6710);
   U4429 : AO4 port map( A => n6655, B => n231, C => n2150, D => n233, Z => 
                           n6711);
   U4430 : AO4 port map( A => n6656, B => n231, C => n2177, D => n233, Z => 
                           n6712);
   U4431 : EOI port map( A => n6657, B => i_SRAM_ADDR_WR05, Z => n2297);
   U4432 : AO4 port map( A => n6658, B => n231, C => i_SRAM_ADDR_WR05, D => 
                           n233, Z => n6714);
   U4433 : AO2 port map( A => KEY_I(0), B => n2430, C => n315, D => 
                           v_KEY32_IN_16_port, Z => n313);
   U4434 : AO2 port map( A => KEY_I(1), B => n2430, C => n315, D => 
                           v_KEY32_IN_17_port, Z => n316);
   U4435 : AO2 port map( A => KEY_I(2), B => n2430, C => n315, D => 
                           v_KEY32_IN_18_port, Z => n317);
   U4436 : AO2 port map( A => KEY_I(3), B => n2430, C => n315, D => 
                           v_KEY32_IN_19_port, Z => n318);
   U4437 : AO2 port map( A => KEY_I(4), B => n2430, C => n315, D => 
                           v_KEY32_IN_20_port, Z => n319);
   U4438 : AO2 port map( A => KEY_I(5), B => n2430, C => n315, D => 
                           v_KEY32_IN_21_port, Z => n320);
   U4439 : AO2 port map( A => KEY_I(6), B => n2430, C => n315, D => 
                           v_KEY32_IN_22_port, Z => n321);
   U4440 : AO2 port map( A => KEY_I(7), B => n2430, C => n315, D => 
                           v_KEY32_IN_23_port, Z => n322);
   U4441 : AO6 port map( A => VALID_KEY_I, B => n4563, C => RESET_I, Z => n239)
                           ;
   U4442 : AO4 port map( A => n2506, B => n333, C => n1832, D => n334, Z => 
                           n6762);
   U4443 : AO6 port map( A => n2505, B => VALID_KEY_I, C => n2391, Z => n333);
   U4444 : AO4 port map( A => n2505, B => CE_I, C => n6803, D => n1719, Z => 
                           n6763);
   U4445 : AO7 port map( A => n4563, B => CE_I, C => n6803, Z => n4604);
   U4446 : IVI port map( A => n707, Z => n2327);
   U4447 : IVI port map( A => n663, Z => n2328);
   U4448 : IVI port map( A => n619, Z => n2329);
   U4449 : IVI port map( A => n575, Z => n2330);
   U4450 : IVI port map( A => n1411, Z => n2331);
   U4451 : IVI port map( A => n1367, Z => n2332);
   U4452 : IVI port map( A => n1323, Z => n2333);
   U4453 : IVI port map( A => n1279, Z => n2334);
   U4454 : IVI port map( A => n531, Z => n2335);
   U4455 : IVI port map( A => n487, Z => n2336);
   U4456 : IVI port map( A => n443, Z => n2337);
   U4457 : IVI port map( A => n442, Z => n2338);
   U4458 : IVI port map( A => n1235, Z => n2339);
   U4459 : IVI port map( A => n1191, Z => n2340);
   U4460 : IVI port map( A => n1147, Z => n2341);
   U4461 : IVI port map( A => n1103, Z => n2342);
   U4462 : IVI port map( A => n441, Z => n2343);
   U4463 : IVI port map( A => n440, Z => n2344);
   U4464 : IVI port map( A => n439, Z => n2345);
   U4465 : IVI port map( A => n438, Z => n2346);
   U4466 : IVI port map( A => n1059, Z => n2347);
   U4467 : IVI port map( A => n1015, Z => n2348);
   U4468 : IVI port map( A => n971, Z => n2349);
   U4469 : IVI port map( A => n927, Z => n2350);
   U4470 : IVI port map( A => n437, Z => n2351);
   U4471 : IVI port map( A => n436, Z => n2352);
   U4472 : IVI port map( A => n435, Z => n2353);
   U4473 : IVI port map( A => n430, Z => n2354);
   U4474 : IVI port map( A => n883, Z => n2355);
   U4475 : IVI port map( A => n839, Z => n2356);
   U4476 : IVI port map( A => n795, Z => n2357);
   U4477 : IVI port map( A => n751, Z => n2358);
   U4478 : IVI port map( A => n429, Z => n2359);
   U4479 : IVI port map( A => n428, Z => n2360);
   U4480 : IVI port map( A => n427, Z => n2361);
   U4481 : IVI port map( A => n426, Z => n2362);
   U4482 : IVI port map( A => n425, Z => n2363);
   U4483 : IVI port map( A => n424, Z => n2364);
   U4484 : IVI port map( A => n423, Z => n2365);
   U4485 : IVI port map( A => n418, Z => n2366);
   U4486 : IVI port map( A => n417, Z => n2367);
   U4488 : IVI port map( A => n416, Z => n2368);
   U4489 : IVI port map( A => n415, Z => n2369);
   U4490 : IVI port map( A => n414, Z => n2370);
   U4491 : IVI port map( A => n413, Z => n2371);
   U4492 : IVI port map( A => n412, Z => n2372);
   U4493 : IVI port map( A => n411, Z => n2373);
   U4494 : IVI port map( A => n406, Z => n2374);
   U4495 : IVI port map( A => n405, Z => n2375);
   U4496 : IVI port map( A => n404, Z => n2376);
   U4497 : IVI port map( A => n403, Z => n2377);
   U4498 : IVI port map( A => n402, Z => n2378);
   U4499 : IVI port map( A => n401, Z => n2379);
   U4500 : IVI port map( A => n400, Z => n2380);
   U4501 : IVI port map( A => n399, Z => n2381);
   U4502 : IVI port map( A => n390, Z => n2382);
   U4503 : IVI port map( A => n389, Z => n2383);
   U4504 : IVI port map( A => n388, Z => n2384);
   U4505 : IVI port map( A => n387, Z => n2385);
   U4506 : IVI port map( A => n386, Z => n2386);
   U4507 : IVI port map( A => n385, Z => n2387);
   U4508 : IVI port map( A => n384, Z => n2388);
   U4509 : IVI port map( A => n383, Z => n2389);
   U4510 : IVI port map( A => n378, Z => n2390);
   U4511 : IVI port map( A => CE_I, Z => n2391);
   U4513 : ND2 port map( A => i_INTERN_ADDR_RD04, B => i_INTERN_ADDR_RD05, Z =>
                           n2392);
   U4514 : AN3 port map( A => i_INTERN_ADDR_RD04, B => i_INTERN_ADDR_RD05, C =>
                           i_INTERN_ADDR_RD03, Z => n2393);
   U4515 : ND2 port map( A => i_INTERN_ADDR_RD02, B => n2393, Z => n2394);
   U4516 : NR2 port map( A => n2394, B => n6660, Z => n2395);
   U4517 : ND2 port map( A => i_SRAM_ADDR_WR04, B => i_SRAM_ADDR_WR05, Z => 
                           n2396);
   U4518 : AN3 port map( A => i_SRAM_ADDR_WR04, B => i_SRAM_ADDR_WR05, C => 
                           i_SRAM_ADDR_WR03, Z => n2397);
   U4519 : ND2 port map( A => i_SRAM_ADDR_WR02, B => n2397, Z => n2398);
   U4520 : NR2 port map( A => n2398, B => n6654, Z => n2399);
   U4521 : ND2 port map( A => v_CALCULATION_CNTR_1_port, B => 
                           v_CALCULATION_CNTR_0_port, Z => n2400);
   U4522 : EN port map( A => v_CALCULATION_CNTR_2_port, B => n2400, Z => N1749)
                           ;
   U4523 : AN3 port map( A => v_CALCULATION_CNTR_1_port, B => 
                           v_CALCULATION_CNTR_0_port, C => 
                           v_CALCULATION_CNTR_2_port, Z => n2402);
   U4524 : EO port map( A => v_CALCULATION_CNTR_3_port, B => n2402, Z => N1750)
                           ;
   U4525 : ND2 port map( A => v_CALCULATION_CNTR_3_port, B => n2402, Z => n2401
                           );
   U4526 : EN port map( A => v_CALCULATION_CNTR_4_port, B => n2401, Z => N1751)
                           ;
   U4527 : AN3 port map( A => v_CALCULATION_CNTR_3_port, B => n2402, C => 
                           v_CALCULATION_CNTR_4_port, Z => n2403);
   U4528 : EO port map( A => v_CALCULATION_CNTR_5_port, B => n2403, Z => N1752)
                           ;
   U4529 : ND2 port map( A => v_CALCULATION_CNTR_5_port, B => n2403, Z => n2404
                           );
   U4530 : EN port map( A => v_CALCULATION_CNTR_6_port, B => n2404, Z => N1753)
                           ;
   U4531 : NR2 port map( A => n2404, B => n2161, Z => n2405);
   U4532 : EO port map( A => v_CALCULATION_CNTR_7_port, B => n2405, Z => N1754)
                           ;
   U4533 : IVI port map( A => n291, Z => n2406);
   U4534 : IVI port map( A => n294, Z => n2407);
   U4535 : IVI port map( A => n295, Z => n2408);
   U4536 : IVI port map( A => n296, Z => n2409);
   U4538 : IVI port map( A => n297, Z => n2410);
   U4539 : IVI port map( A => n298, Z => n2411);
   U4540 : IVI port map( A => n299, Z => n2412);
   U4541 : IVI port map( A => n300, Z => n2413);
   U4542 : IVI port map( A => n323, Z => n2414);
   U4543 : IVI port map( A => n326, Z => n2415);
   U4544 : IVI port map( A => n327, Z => n2416);
   U4545 : IVI port map( A => n328, Z => n2417);
   U4546 : IVI port map( A => n329, Z => n2418);
   U4547 : IVI port map( A => n330, Z => n2419);
   U4548 : IVI port map( A => n331, Z => n2420);
   U4549 : IVI port map( A => n332, Z => n2421);
   U4550 : IVI port map( A => n313, Z => n2422);
   U4551 : IVI port map( A => n316, Z => n2423);
   U4552 : IVI port map( A => n317, Z => n2424);
   U4553 : IVI port map( A => n318, Z => n2425);
   U4554 : IVI port map( A => n319, Z => n2426);
   U4555 : IVI port map( A => n320, Z => n2427);
   U4556 : IVI port map( A => n321, Z => n2428);
   U4557 : IVI port map( A => n322, Z => n2429);
   U4558 : IVI port map( A => n315, Z => n2430);
   U4559 : IVI port map( A => n302, Z => n2431);
   U4560 : IVI port map( A => n305, Z => n2432);
   U4561 : IVI port map( A => n306, Z => n2433);
   U4563 : IVI port map( A => n307, Z => n2434);
   U4564 : IVI port map( A => n308, Z => n2435);
   U4565 : IVI port map( A => n309, Z => n2436);
   U4567 : IVI port map( A => n310, Z => n2437);
   U4568 : IVI port map( A => n311, Z => n2438);
   U4569 : IVI port map( A => n279, Z => n2479);
   U4571 : IVI port map( A => n268, Z => n2481);
   U4572 : IVI port map( A => n2500, Z => n2491);
   U4573 : IVI port map( A => n2502, Z => n2492);
   U4575 : IVI port map( A => n2503, Z => n2494);
   U4576 : IVI port map( A => n57, Z => n2501);
   U4577 : IVI port map( A => n64, Z => n2504);
   U4579 : IVI port map( A => n1951, Z => n2508);
   U4580 : IVI port map( A => n1850, Z => n4558);
   U4581 : IVI port map( A => n1953, Z => n4559);
   U4582 : IVI port map( A => n2026, Z => n4560);
   U4583 : IVI port map( A => n2119, Z => n4562);
   U4584 : IVI port map( A => n2128, Z => n6670);
   U4585 : IVI port map( A => n2182, Z => n6671);
   U4586 : IVI port map( A => n2151, Z => n6672);
   U4587 : IVI port map( A => n2011, Z => n6730);
   U4588 : IVI port map( A => n2058, Z => n6731);
   U4589 : IVI port map( A => n2239, Z => n6732);
   U4590 : IVI port map( A => n2028, Z => n6734);
   U4591 : IVI port map( A => n2118, Z => n6735);
   U4592 : IVI port map( A => n1971, Z => n6736);
   U4593 : IVI port map( A => n2032, Z => n6737);
   U4594 : IVI port map( A => n2129, Z => n6738);
   U4595 : IVI port map( A => n1940, Z => n6739);
   U4597 : IVI port map( A => n1939, Z => n6740);
   U4601 : IVI port map( A => n1930, Z => n6741);
   U4605 : IVI port map( A => n2282, Z => n6742);
   U4606 : IVI port map( A => n2162, Z => n6743);
   U4607 : IVI port map( A => n2208, Z => n6744);
   U4608 : IVI port map( A => n2002, Z => n6745);
   U4609 : IVI port map( A => n1909, Z => n6746);
   U4610 : IVI port map( A => n2049, Z => n6748);
   U4611 : IVI port map( A => n2188, Z => n6749);
   U4614 : IVI port map( A => n2246, Z => n6750);
   U4616 : IVI port map( A => n1859, Z => n6751);
   U4617 : IVI port map( A => n1988, Z => n6752);
   U4618 : IVI port map( A => n2010, Z => n6753);
   U4619 : IVI port map( A => n1887, Z => n6754);
   U4620 : IVI port map( A => n1969, Z => n6755);
   U4621 : IVI port map( A => n2043, Z => n6756);
   U4622 : IVI port map( A => n1944, Z => n6757);
   U4623 : IVI port map( A => n1895, Z => n6758);
   U4624 : IVI port map( A => n2084, Z => n6759);
   U4625 : IVI port map( A => n2187, Z => n6760);
   U4626 : IVI port map( A => n2178, Z => n6761);
   U4627 : IVI port map( A => n2051, Z => n6765);
   U4628 : IVI port map( A => n2000, Z => n6766);
   U4629 : IVI port map( A => n2102, Z => n6767);
   U4630 : IVI port map( A => n1885, Z => n6768);
   U4631 : IVI port map( A => n1938, Z => n6769);
   U4632 : IVI port map( A => n2039, Z => n6770);
   U4633 : IVI port map( A => n2093, Z => n6771);
   U4634 : IVI port map( A => n2024, Z => n6772);
   U4636 : IVI port map( A => n1998, Z => n6773);
   U4637 : IVI port map( A => n1886, Z => n6775);
   U4638 : IVI port map( A => n1897, Z => n6777);
   U4640 : IVI port map( A => n2105, Z => n6778);
   U4641 : IVI port map( A => n2184, Z => n6779);
   U4643 : IVI port map( A => n1980, Z => n6780);
   U4644 : IVI port map( A => n149, Z => n6781);
   U4646 : IVI port map( A => n154, Z => n6782);
   U4648 : IVI port map( A => n108, Z => n6783);
   U4650 : IVI port map( A => n113, Z => n6784);
   U4652 : IVI port map( A => n171, Z => n6785);
   U4654 : IVI port map( A => n267, Z => n6786);
   U4656 : IVI port map( A => n290, Z => n6787);
   U4658 : IVI port map( A => n282, Z => n6788);
   U4660 : IVI port map( A => n2299, Z => n6789);
   U4662 : IVI port map( A => n155, Z => n6790);
   U4664 : IVI port map( A => n65, Z => n6791);
   U4666 : IVI port map( A => n169, Z => n6792);
   U4668 : IVI port map( A => n2307, Z => n6793);
   U4670 : IVI port map( A => n266, Z => n6794);
   U4672 : IVI port map( A => n2498, Z => n6795);
   U4674 : IVI port map( A => n1845, Z => n6796);
   U4676 : IVI port map( A => n1846, Z => n6797);
   U4678 : IVI port map( A => n1835, Z => n6798);
   U4680 : IVI port map( A => n1836, Z => n6799);
   U4682 : IVI port map( A => n1807, Z => n6800);
   U4684 : IVI port map( A => n1808, Z => n6801);
   U4686 : IVI port map( A => n2485, Z => n6802);
   U4688 : IVI port map( A => n263, Z => n6803);
   U4690 : IVI port map( A => VALID_KEY_I, Z => n6804);
   U4692 : IVI port map( A => n242, Z => n6805);
   U4694 : IVI port map( A => RESET_I, Z => n6806);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_aes_dec_KEY_SIZE2.all;

entity aes_dec_KEY_SIZE2 is

   port( DATA_I : in std_logic_vector (7 downto 0);  VALID_DATA_I : in 
         std_logic;  KEY_I : in std_logic_vector (7 downto 0);  VALID_KEY_I, 
         RESET_I, CLK_I, CE_I : in std_logic;  KEY_READY_O, VALID_O : out 
         std_logic;  DATA_O : out std_logic_vector (7 downto 0));

end aes_dec_KEY_SIZE2;

architecture SYN_Behavioral of aes_dec_KEY_SIZE2 is

   component IVI
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component EO
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NR2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EN
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component ND2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AN3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component AO7
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component IV
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AO6
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component IVA
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AO4
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component EON1
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component AO2
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component AO3
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component IVDA
      port( A : in std_logic;  Y, Z : out std_logic);
   end component;
   
   component ND4
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component NR3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component ND2I
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EOI
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NR4
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component EO1
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component ND3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component ENI
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AN2I
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NR2I
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component key_expansion
      port( KEY_I : in std_logic_vector (7 downto 0);  VALID_KEY_I, CLK_I, 
            RESET_I, CE_I : in std_logic;  DONE_O : out std_logic;  GET_KEY_I :
            in std_logic;  KEY_NUMB_I : in std_logic_vector (5 downto 0);  
            KEY_EXP_O : out std_logic_vector (31 downto 0));
   end component;
   
   component AO1P
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OR4
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component FD1
      port( D, CP : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal DATA_O_7_port, DATA_O_6_port, DATA_O_5_port, DATA_O_4_port, 
      DATA_O_3_port, DATA_O_2_port, DATA_O_1_port, DATA_O_0_port, GET_KEY, 
      v_INV_KEY_NUMB_5_port, v_INV_KEY_NUMB_4_port, v_INV_KEY_NUMB_3_port, 
      v_INV_KEY_NUMB_2_port, v_KEY_COLUMN_31_port, v_KEY_COLUMN_30_port, 
      v_KEY_COLUMN_29_port, v_KEY_COLUMN_28_port, v_KEY_COLUMN_27_port, 
      v_KEY_COLUMN_26_port, v_KEY_COLUMN_25_port, v_KEY_COLUMN_24_port, 
      v_KEY_COLUMN_23_port, v_KEY_COLUMN_22_port, v_KEY_COLUMN_21_port, 
      v_KEY_COLUMN_20_port, v_KEY_COLUMN_19_port, v_KEY_COLUMN_18_port, 
      v_KEY_COLUMN_17_port, v_KEY_COLUMN_16_port, v_KEY_COLUMN_15_port, 
      v_KEY_COLUMN_14_port, v_KEY_COLUMN_13_port, v_KEY_COLUMN_12_port, 
      v_KEY_COLUMN_11_port, v_KEY_COLUMN_10_port, v_KEY_COLUMN_9_port, 
      v_KEY_COLUMN_8_port, v_KEY_COLUMN_7_port, v_KEY_COLUMN_6_port, 
      v_KEY_COLUMN_5_port, v_KEY_COLUMN_4_port, v_KEY_COLUMN_3_port, 
      v_KEY_COLUMN_2_port, v_KEY_COLUMN_1_port, v_KEY_COLUMN_0_port, 
      v_CNT4_1_port, v_CNT4_0_port, v_DATA_COLUMN_31_port, 
      v_DATA_COLUMN_30_port, v_DATA_COLUMN_29_port, v_DATA_COLUMN_28_port, 
      v_DATA_COLUMN_27_port, v_DATA_COLUMN_26_port, v_DATA_COLUMN_25_port, 
      v_DATA_COLUMN_24_port, v_DATA_COLUMN_23_port, v_DATA_COLUMN_22_port, 
      v_DATA_COLUMN_21_port, v_DATA_COLUMN_20_port, v_DATA_COLUMN_19_port, 
      v_DATA_COLUMN_18_port, v_DATA_COLUMN_17_port, v_DATA_COLUMN_16_port, 
      v_DATA_COLUMN_15_port, v_DATA_COLUMN_14_port, v_DATA_COLUMN_13_port, 
      v_DATA_COLUMN_12_port, v_DATA_COLUMN_11_port, v_DATA_COLUMN_10_port, 
      v_DATA_COLUMN_9_port, v_DATA_COLUMN_8_port, v_DATA_COLUMN_7_port, 
      v_DATA_COLUMN_6_port, v_DATA_COLUMN_5_port, v_DATA_COLUMN_4_port, 
      v_DATA_COLUMN_3_port, v_DATA_COLUMN_2_port, v_DATA_COLUMN_1_port, 
      v_DATA_COLUMN_0_port, v_CALCULATION_CNTR_7_port, 
      v_CALCULATION_CNTR_6_port, v_CALCULATION_CNTR_5_port, 
      v_CALCULATION_CNTR_4_port, v_CALCULATION_CNTR_3_port, 
      v_CALCULATION_CNTR_2_port, v_CALCULATION_CNTR_1_port, 
      v_CALCULATION_CNTR_0_port, N192, N199, N200, N201, N202, N203, 
      t_STATE_RAM0_0_31_port, t_STATE_RAM0_0_30_port, t_STATE_RAM0_0_29_port, 
      t_STATE_RAM0_0_28_port, t_STATE_RAM0_0_27_port, t_STATE_RAM0_0_26_port, 
      t_STATE_RAM0_0_25_port, t_STATE_RAM0_0_24_port, t_STATE_RAM0_0_23_port, 
      t_STATE_RAM0_0_22_port, t_STATE_RAM0_0_21_port, t_STATE_RAM0_0_20_port, 
      t_STATE_RAM0_0_19_port, t_STATE_RAM0_0_18_port, t_STATE_RAM0_0_17_port, 
      t_STATE_RAM0_0_16_port, t_STATE_RAM0_0_15_port, t_STATE_RAM0_0_14_port, 
      t_STATE_RAM0_0_13_port, t_STATE_RAM0_0_12_port, t_STATE_RAM0_0_11_port, 
      t_STATE_RAM0_0_10_port, t_STATE_RAM0_0_9_port, t_STATE_RAM0_0_8_port, 
      t_STATE_RAM0_0_7_port, t_STATE_RAM0_0_6_port, t_STATE_RAM0_0_5_port, 
      t_STATE_RAM0_0_4_port, t_STATE_RAM0_0_3_port, t_STATE_RAM0_0_2_port, 
      t_STATE_RAM0_0_1_port, t_STATE_RAM0_0_0_port, t_STATE_RAM0_1_31_port, 
      t_STATE_RAM0_1_30_port, t_STATE_RAM0_1_29_port, t_STATE_RAM0_1_28_port, 
      t_STATE_RAM0_1_27_port, t_STATE_RAM0_1_26_port, t_STATE_RAM0_1_25_port, 
      t_STATE_RAM0_1_24_port, t_STATE_RAM0_1_23_port, t_STATE_RAM0_1_22_port, 
      t_STATE_RAM0_1_21_port, t_STATE_RAM0_1_20_port, t_STATE_RAM0_1_19_port, 
      t_STATE_RAM0_1_18_port, t_STATE_RAM0_1_17_port, t_STATE_RAM0_1_16_port, 
      t_STATE_RAM0_1_15_port, t_STATE_RAM0_1_14_port, t_STATE_RAM0_1_13_port, 
      t_STATE_RAM0_1_12_port, t_STATE_RAM0_1_11_port, t_STATE_RAM0_1_10_port, 
      t_STATE_RAM0_1_9_port, t_STATE_RAM0_1_8_port, t_STATE_RAM0_1_7_port, 
      t_STATE_RAM0_1_6_port, t_STATE_RAM0_1_5_port, t_STATE_RAM0_1_4_port, 
      t_STATE_RAM0_1_3_port, t_STATE_RAM0_1_2_port, t_STATE_RAM0_1_1_port, 
      t_STATE_RAM0_1_0_port, t_STATE_RAM0_2_31_port, t_STATE_RAM0_2_30_port, 
      t_STATE_RAM0_2_29_port, t_STATE_RAM0_2_28_port, t_STATE_RAM0_2_27_port, 
      t_STATE_RAM0_2_26_port, t_STATE_RAM0_2_25_port, t_STATE_RAM0_2_24_port, 
      t_STATE_RAM0_2_23_port, t_STATE_RAM0_2_22_port, t_STATE_RAM0_2_21_port, 
      t_STATE_RAM0_2_20_port, t_STATE_RAM0_2_19_port, t_STATE_RAM0_2_18_port, 
      t_STATE_RAM0_2_17_port, t_STATE_RAM0_2_16_port, t_STATE_RAM0_2_15_port, 
      t_STATE_RAM0_2_14_port, t_STATE_RAM0_2_13_port, t_STATE_RAM0_2_12_port, 
      t_STATE_RAM0_2_11_port, t_STATE_RAM0_2_10_port, t_STATE_RAM0_2_9_port, 
      t_STATE_RAM0_2_8_port, t_STATE_RAM0_2_7_port, t_STATE_RAM0_2_6_port, 
      t_STATE_RAM0_2_5_port, t_STATE_RAM0_2_4_port, t_STATE_RAM0_2_3_port, 
      t_STATE_RAM0_2_2_port, t_STATE_RAM0_2_1_port, t_STATE_RAM0_2_0_port, 
      v_RAM_OUT0_31_port, v_RAM_OUT0_30_port, v_RAM_OUT0_29_port, 
      v_RAM_OUT0_28_port, v_RAM_OUT0_27_port, v_RAM_OUT0_26_port, 
      v_RAM_OUT0_25_port, v_RAM_OUT0_24_port, v_RAM_OUT0_23_port, 
      v_RAM_OUT0_22_port, v_RAM_OUT0_21_port, v_RAM_OUT0_20_port, 
      v_RAM_OUT0_19_port, v_RAM_OUT0_18_port, v_RAM_OUT0_17_port, 
      v_RAM_OUT0_16_port, v_RAM_OUT0_15_port, v_RAM_OUT0_14_port, 
      v_RAM_OUT0_13_port, v_RAM_OUT0_12_port, v_RAM_OUT0_11_port, 
      v_RAM_OUT0_10_port, v_RAM_OUT0_9_port, v_RAM_OUT0_8_port, 
      v_RAM_OUT0_7_port, v_RAM_OUT0_6_port, v_RAM_OUT0_5_port, 
      v_RAM_OUT0_4_port, v_RAM_OUT0_3_port, v_RAM_OUT0_2_port, 
      v_RAM_OUT0_1_port, v_RAM_OUT0_0_port, N2083, N2084, N2085, N2086, N2087, 
      N2088, N2089, n3, n4, n10, n11, n13, n14, n16, n17, n19, n20, n22, n23, 
      n25, n26, n28, n29, n31, n32, n34, n35, n37, n38, n40, n41, n43, n44, n46
      , n47, n49, n50, n52, n53, n55, n56, n58, n59, n61, n62, n64, n65, n67, 
      n68, n70, n71, n73, n74, n76, n77, n79, n80, n82, n83, n85, n86, n88, n89
      , n91, n92, n94, n95, n97, n98, n100, n101, n103, n105, n107, n108, n109,
      n111, n113, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, 
      n125, n126, n127, n128, n129, n130, n131, n132, n133, n135, n136, n138, 
      n139, n140, n141, n142, n143, n145, n146, n147, n149, n150, n151, n152, 
      n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n164, n165, 
      n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n177, n178, 
      n179, n180, n181, n182, n183, n184, n185, n186, n188, n189, n190, 
      n192_port, n195, n196, n197, n199_port, n201_port, n202_port, n203_port, 
      n204, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, 
      n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, 
      n229, n230, n231, n232, n233, n235, n236, n237, n238, n239, n240, n241, 
      n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, 
      n254, n255, n256, n257, n258, n260, n261, n262, n263, n264, n265, n266, 
      n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
      n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
      n291, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, 
      n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, 
      n316, n317, n318, n319, n320, n321, n322, n323, n324, n326, n327, n328, 
      n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, 
      n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, 
      n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, 
      n365, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, 
      n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, 
      n390, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n425, n426, n427, 
      n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, 
      n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, 
      n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, 
      n464, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, 
      n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, 
      n489, n490, n491, n492, n493, n494, n495, n496, n497, n499, n500, n501, 
      n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, 
      n514, n515, n516, n517, n518, n519, n520, n521, n522, n524, n525, n526, 
      n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, 
      n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n551, 
      n552, n553, n554, n555, n556, n557, n558, n559, n561, n563, n564, n565, 
      n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, 
      n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, 
      n590, n591, n592, n593, n594, n596, n597, n598, n599, n600, n601, n602, 
      n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n614, n615, 
      n616, n617, n618, n621, n622, n623, n624, n625, n626, n627, n628, n629, 
      n630, n631, n632, n633, n634, n635, n636, n638, n639, n640, n641, n642, 
      n643, n644, n645, n646, n647, n648, n649, n650, n652, n653, n654, n655, 
      n656, n657, n658, n659, n660, n661, n664, n665, n666, n667, n668, n669, 
      n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, 
      n682, n683, n684, n686, n687, n688, n689, n691, n692, n693, n694, n695, 
      n696, n697, n700, n702, n703, n704, n705, n706, n707, n708, n709, n710, 
      n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, 
      n723, n724, n725, n726, n727, n728, n729, n731, n732, n733, n734, n735, 
      n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, 
      n748, n749, n750, n751, n752, n753, n754, n756, n757, n758, n759, n760, 
      n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, 
      n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, 
      n785, n786, n787, n788, n789, n790, n793, n794, n795, n796, n797, n798, 
      n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, 
      n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, 
      n823, n824, n825, n826, n827, n828, n829, n831, n832, n833, n835, n836, 
      n837, n838, n839, n840, n841, n842, n843, n844, n846, n847, n848, n849, 
      n850, n851, n852, n853, n854, n855, n857, n858, n859, n860, n861, n862, 
      n863, n864, n865, n866, n867, n868, n869, n870, n871, n873, n874, n875, 
      n876, n877, n878, n879, n880, n881, n882, n883, n884, n886, n888, n889, 
      n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, 
      n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, 
      n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, 
      n926, n928, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, 
      n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, 
      n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n964, 
      n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, 
      n978, n979, n980, n981, n982, n983, n984, n985, n987, n988, n989, n990, 
      n991, n992, n994, n995, n996, n998, n1001, n1003, n1004, n1007, n1008, 
      n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1017, n1018, n1019, 
      n1022, n1023, n1024, n1027, n1028, n1029, n1030, n1031, n1033, n1036, 
      n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1046, n1047, 
      n1048, n1049, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, 
      n1059, n1060, n1061, n1062, n1063, n1065, n1066, n1067, n1068, n1069, 
      n1070, n1071, n1072, n1073, n1075, n1076, n1079, n1080, n1081, n1083, 
      n1084, n1086, n1087, n1088, n1090, n1092, n1093, n1094, n1095, n1096, 
      n1097, n1100, n1101, n1102, n1104, n1105, n1106, n1107, n1108, n1109, 
      n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1119, n1122, n1124, 
      n1125, n1126, n1127, n1128, n1129, n1130, n1132, n1134, n1136, n1137, 
      n1139, n1140, n1141, n1142, n1143, n1145, n1147, n1148, n1149, n1150, 
      n1151, n1153, n1154, n1155, n1156, n1157, n1160, n1162, n1164, n1165, 
      n1166, n1167, n1168, n1169, n1170, n1171, n1175, n1176, n1177, n1178, 
      n1185, n1189, n1190, n1193, n1194, n1195, n1196, n1203, n1206, n1207, 
      n1208, n1211, n1212, n1213, n1214, n1221, n1222, n1223, n1224, n1225, 
      n1229, n1230, n1231, n1232, n1240, n1241, n1242, n1243, n1245, n1246, 
      n1247, n1251, n1252, n1253, n1254, n1257, n1265, n1266, n1269, n1270, 
      n1271, n1272, n1275, n1280, n1281, n1282, n1283, n1284, n1287, n1289, 
      n1293, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1306, n1307, 
      n1313, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1339, 
      n1340, n1341, n1342, n1350, n1351, n1353, n1354, n1355, n1356, n1364, 
      n1365, n1366, n1370, n1371, n1374, n1376, n1386, n1387, n1391, n1392, 
      n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1403, n1404, 
      n1406, n1407, n1408, n1410, n1411, n1412, n1413, n1414, n1415, n1417, 
      n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, 
      n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, 
      n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1447, n1448, n1450, 
      n1451, n1452, n1454, n1459, n1465, n1467, n1469, n1470, n1471, n1474, 
      n1475, n1476, n1477, n1480, n1481, n1482, n1483, n1485, n1486, n1487, 
      n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1498, n1499, n1501, 
      n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, 
      n1513, n1515, n1516, n1517, n1520, n1521, n1522, n1523, n1524, n1525, 
      n1527, n1528, n1529, n1530, n1531, n1532, n1534, n1535, n1536, n1537, 
      n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1548, n1549, 
      n1550, n1551, n1552, n1553, n1554, n1555, n1557, n1558, n1559, n1560, 
      n1561, n1562, n1563, n1564, n1565, n1566, n1568, n1569, n1570, n1571, 
      n1572, n1574, n1576, n1577, n1580, n1581, n1582, n1583, n1584, n1585, 
      n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, 
      n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, 
      n1609, n1610, n1611, n1612, n1613, n1614, n1616, n1618, n1619, n1620, 
      n1621, n1622, n1623, n1626, n1627, n1628, n1629, n1631, n1632, n1633, 
      n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1644, 
      n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1656, 
      n1658, n1659, n1660, n1661, n1662, n1663, n1666, n1667, n1668, n1669, 
      n1670, n1671, n1672, n1673, n1674, n1675, n1679, n1680, n1684, n1685, 
      n1686, n1687, n1688, n1689, n1694, n1695, n1696, n1697, n1698, n1699, 
      n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1710, n1711, 
      n1712, n1713, n1716, n1717, n1719, n1720, n1722, n1723, n1724, n1725, 
      n1726, n1727, n1728, n1730, n1731, n1732, n1733, n1734, n1735, n1736, 
      n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, 
      n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, 
      n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1766, n1767, n1768, 
      n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1779, 
      n1780, n1781, n1782, n1783, n1784, n1785, n1787, n1788, n1789, n1790, 
      n1791, n1792, n1793, n1794, n1795, n1796, n1798, n1799, n1800, n1801, 
      n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, 
      n1812, n1813, n1814, n1815, n1816, n1817, n1819, n1820, n1821, n1822, 
      n1823, n1824, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, 
      n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, 
      n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1853, n1854, n1855, 
      n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1865, n1866, 
      n1867, n1868, n1869, n1870, n1872, n1876, n1877, n1878, n1879, n1882, 
      n1883, n1885, n1886, n1887, n1888, n1889, n1890, n1892, n1893, n1894, 
      n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1904, n1906, 
      n1907, n1909, n1910, n1911, n1912, n1913, n1914, n1916, n1917, n1918, 
      n1919, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1930, n1931, 
      n1932, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1942, n1944, 
      n1945, n1947, n1948, n1949, n1951, n1952, n1953, n1955, n1958, n1959, 
      n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, 
      n1970, n1973, n1974, n1975, n1977, n1978, n1980, n1982, n1983, n1985, 
      n1986, n1987, n1988, n1991, n1992, n1993, n1994, n1995, n1997, n1999, 
      n2002, n2003, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, 
      n2013, n2014, n2015, n2016, n2017, n2019, n2020, n2021, n2022, n2023, 
      n2024, n2025, n2026, n2027, n2028, n2029, n2031, n2032, n2033, n2035, 
      n2038, n2040, n2041, n2043, n2044, n2046, n2047, n2048, n2050, n2051, 
      n2052, n2054, n2055, n2056, n2057, n2058, n2060, n2061, n2064, n2065, 
      n2066, n2067, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, 
      n2077, n2082, n2083_port, n2084_port, n2085_port, n2087_port, n2089_port,
      n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2101, 
      n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, 
      n2112, n2113, n2114, n2117, n2118, n2119, n2120, n2121, n2123, n2124, 
      n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2133, n2136, n2137, 
      n2138, n2139, n2140, n2141, n2142, n2144, n2145, n2146, n2147, n2148, 
      n2150, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2162, 
      n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, 
      n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, 
      n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, 
      n2194, n2195, n2196, n2197, n2198, n2199, n2201, n2202, n2203, n2204, 
      n2205, n2206, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, 
      n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, 
      n2227, n2228, n2230, n2231, n2232, n2233, n2234, n2236, n2237, n2238, 
      n2239, n2241, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, 
      n2251, n2252, n2253, n2256, n2257, n2259, n2260, n2261, n2262, n2264, 
      n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2274, n2275, 
      n2276, n2277, n2278, n2279, n2281, n2282, n2283, n2285, n2286, n2287, 
      n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2296, n2297, n2298, 
      n2299, n2300, n2301, n2302, n2304, n2305, n2306, n2307, n2308, n2309, 
      n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, 
      n2321, n2322, n2323, n2324, n2325, n2327, n2328, n2329, n2330, n2331, 
      n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, 
      n2342, n2343, n2344, n2345, n2346, n2347, n2349, n2350, n2351, n2352, 
      n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, 
      n2363, n2364, n2365, n2367, n2369, n2370, n2372, n2373, n2374, n2375, 
      n2376, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, 
      n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, 
      n2397, n2398, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, 
      n2410, n2411, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, 
      n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, 
      n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, 
      n2441, n2445, n2446, n2450, n2451, n2452, n2453, n2454, n2455, n2460, 
      n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, 
      n2471, n2474, n2475, n2476, n2477, n2480, n2481, n2483, n2484, n2486, 
      n2487, n2488, n2489, n2490, n2491, n2492, n2494, n2495, n2496, n2497, 
      n2498, n2499, n2500, n2501, n2502, n2503, n2505, n2507, n2509, n2510, 
      n2513, n2515, n2516, n2517, n2519, n2520, n2521, n2522, n2523, n2525, 
      n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2536, n2537, 
      n2538, n2539, n2540, n2541, n2542, n2544, n2547, n2548, n2549, n2550, 
      n2552, n2553, n2554, n2555, n2557, n2559, n2560, n2561, n2562, n2565, 
      n2567, n2568, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, 
      n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, 
      n2589, n2590, n2591, n2593, n2594, n2595, n2596, n2597, n2598, n2600, 
      n2601, n2605, n2606, n2608, n2609, n2610, n2612, n2615, n2616, n2617, 
      n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, 
      n2628, n2629, n2630, n2632, n2633, n2634, n2635, n2636, n2637, n2638, 
      n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2647, n2648, n2649, 
      n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, 
      n2661, n2662, n2663, n2665, n2666, n2667, n2670, n2672, n2673, n2674, 
      n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, 
      n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2695, n2696, n2698, 
      n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, 
      n2709, n2710, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, 
      n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, 
      n2730, n2731, n2732, n2734, n2735, n2736, n2737, n2738, n2739, n2740, 
      n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, 
      n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, 
      n2761, n2762, n2763, n2764, n2765, n2767, n2768, n2769, n2770, n2771, 
      n2772, n2773, n2774, n2776, n2777, n2778, n2779, n2781, n2782, n2783, 
      n2784, n2785, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, 
      n2795, n2796, n2797, n2798, n2799, n2801, n2802, n2803, n2804, n2805, 
      n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, 
      n2817, n2818, n2819, n2820, n2821, n2822, n2824, n2825, n2826, n2827, 
      n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, 
      n2838, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, 
      n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, 
      n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, 
      n2870, n2871, n2872, n2873, n2874, n2876, n2878, n2879, n2880, n2881, 
      n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, 
      n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, 
      n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2911, n2913, n2914, 
      n2917, n2919, n2920, n2921, n2923, n2924, n2925, n2926, n2927, n2930, 
      n2932, n2933, n2935, n2936, n2938, n2939, n2940, n2942, n2943, n2944, 
      n2945, n2946, n2947, n2949, n2951, n2952, n2953, n2954, n2955, n2956, 
      n2957, n2958, n2959, n2961, n2962, n2963, n2964, n2965, n2968, n2969, 
      n2970, n2971, n2972, n2974, n2975, n2976, n2977, n2978, n2979, n2981, 
      n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2992, 
      n2993, n2995, n2996, n2997, n2998, n2999, n3000, n3002, n3003, n3007, 
      n3008, n3009, n3011, n3012, n3013, n3014, n3017, n3018, n3019, n3020, 
      n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3030, n3031, n3032, 
      n3033, n3034, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, 
      n3044, n3045, n3046, n3047, n3048, n3049, n3051, n3052, n3053, n3055, 
      n3056, n3057, n3058, n3060, n3061, n3062, n3063, n3064, n3065, n3066, 
      n3067, n3068, n3070, n3071, n3072, n3075, n3077, n3078, n3079, n3080, 
      n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3091, 
      n3092, n3093, n3094, n3095, n3096, n3097, n3100, n3101, n3103, n3104, 
      n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, 
      n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, 
      n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, 
      n3135, n3136, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, 
      n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, 
      n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, 
      n3166, n3167, n3168, n3169, n3171, n3172, n3173, n3174, n3175, n3176, 
      n3177, n3178, n3180, n3181, n3182, n3183, n3184, n3186, n3187, n3188, 
      n3189, n3190, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, 
      n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3210, 
      n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3219, n3220, n3221, 
      n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, 
      n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, 
      n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3254, 
      n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, 
      n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, 
      n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3285, 
      n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, 
      n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, 
      n3306, n3307, n3308, n3309, n3310, n3313, n3315, n3316, n3319, n3321, 
      n3322, n3323, n3325, n3326, n3327, n3328, n3329, n3332, n3334, n3335, 
      n3337, n3338, n3340, n3341, n3342, n3344, n3345, n3346, n3347, n3348, 
      n3349, n3351, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, 
      n3361, n3363, n3364, n3365, n3366, n3367, n3370, n3371, n3372, n3373, 
      n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3382, n3383, n3384, 
      n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3393, n3394, n3396, 
      n3397, n3398, n3399, n3400, n3401, n3403, n3404, n3408, n3409, n3410, 
      n3412, n3413, n3414, n3415, n3418, n3419, n3420, n3421, n3423, n3424, 
      n3425, n3426, n3427, n3428, n3429, n3431, n3432, n3433, n3434, n3435, 
      n3437, n3438, n3439, n3440, n3441, n3442, n3444, n3445, n3446, n3447, 
      n3448, n3449, n3450, n3451, n3453, n3454, n3455, n3457, n3458, n3459, 
      n3460, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, 
      n3472, n3473, n3474, n3477, n3479, n3480, n3481, n3482, n3483, n3484, 
      n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3493, n3494, n3495, 
      n3496, n3497, n3498, n3499, n3502, n3503, n3504, n3505, n3506, n3507, 
      n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, 
      n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, 
      n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, 
      n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, 
      n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, 
      n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, 
      n3569, n3570, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, 
      n3581, n3582, n3583, n3584, n3585, n3587, n3588, n3589, n3590, n3591, 
      n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, 
      n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3611, n3612, n3613, 
      n3614, n3615, n3616, n3617, n3618, n3620, n3621, n3622, n3624, n3625, 
      n3626, n3627, n3628, n3629, n3630, n3632, n3633, n3634, n3635, n3636, 
      n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3646, n3647, 
      n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3656, n3657, n3658, 
      n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, 
      n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, 
      n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3689, 
      n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, 
      n3700, n3701, n3703, n3704, n3705, n3706, n3708, n3710, n3712, n3713, 
      n3714, n3715, n3716, n3717, n3718, n3719, n3721, n3722, n3723, n3724, 
      n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, 
      n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, 
      n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, 
      n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, 
      n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, 
      n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, 
      n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, 
      n3795, n3796, n3798, n3799, n3800, n3801, n3802, n3803, n3805, n3806, 
      n3807, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, 
      n3818, n3823, n3824, n3825, n3835, n3836, n3837, n3838, n3839, n3840, 
      n3841, n3842, n3847, n3850, n3851, n3852, n3853, n3854, n3855, n3856, 
      n3857, n3858, n3860, n3864, n3866, n3868, n3872, n3879, n3882, n3887, 
      n3889, n3896, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, 
      n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, 
      n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3924, n3928, n3930, 
      n3932, n3936, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, 
      n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, 
      n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, 
      n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, 
      n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, 
      n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, 
      n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, 
      n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, 
      n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, 
      n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, 
      n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, 
      n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, 
      n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, 
      n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, 
      n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, 
      n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, 
      n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, 
      n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, 
      n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, 
      n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, 
      n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, 
      n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, 
      n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, 
      n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, 
      n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, 
      n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, 
      n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, 
      n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, 
      n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, 
      n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, 
      n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, 
      n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, 
      n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, 
      n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, 
      n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, 
      n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, 
      n4297, n4298, n4300, n4301, n4302, n4306, n4307, n4308, n4309, n4310, 
      n4311, n4312, n4337, n4346, n4349, n4350, n4351, n4352, n4353, n4354, 
      n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, 
      n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, 
      n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, 
      n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, 
      n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, 
      n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, 
      n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, 
      n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, 
      n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, 
      n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, 
      n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, 
      n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, 
      n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, 
      n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, 
      n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, 
      n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, 
      n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, 
      n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, 
      n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, 
      n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, 
      n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, 
      n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, 
      n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, 
      n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, 
      n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, 
      n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, 
      n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, 
      n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, 
      n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, 
      n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, 
      n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, 
      n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, 
      n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, 
      n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, 
      n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, 
      n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, 
      n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, 
      n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, 
      n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, 
      n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, 
      n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, 
      n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, 
      n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, 
      n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, 
      n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, 
      n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, 
      n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, 
      n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, 
      n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, 
      n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, 
      n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, 
      n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, 
      n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, 
      n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, 
      n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, 
      n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, 
      n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, 
      n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, 
      n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, 
      n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, 
      n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, 
      n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, 
      n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, 
      n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, 
      n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, 
      n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, 
      n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, 
      n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, 
      n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, 
      n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, 
      n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, 
      n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n_3156, 
      n_3157, n_3158, n_3159, n_3160, n_3161, n_3162, n_3163, n_3164, n_3165, 
      n_3166, n_3167, n_3168, n_3169, n_3170, n_3171, n_3172, n_3173, n_3174, 
      n_3175, n_3176, n_3177, n_3178, n_3179, n_3180, n_3181, n_3182, n_3183, 
      n_3184, n_3185, n_3186, n_3187, n_3188, n_3189, n_3190, n_3191, n_3192, 
      n_3193, n_3194, n_3195, n_3196, n_3197, n_3198, n_3199, n_3200, n_3201, 
      n_3202, n_3203, n_3204, n_3205, n_3206, n_3207, n_3208, n_3209, n_3210, 
      n_3211, n_3212, n_3213, n_3214, n_3215, n_3216, n_3217, n_3218, n_3219, 
      n_3220, n_3221, n_3222, n_3223, n_3224, n_3225, n_3226, n_3227, n_3228, 
      n_3229, n_3230, n_3231, n_3232, n_3233, n_3234, n_3235, n_3236, n_3237, 
      n_3238, n_3239, n_3240, n_3241, n_3242, n_3243, n_3244, n_3245, n_3246, 
      n_3247, n_3248, n_3249, n_3250, n_3251, n_3252, n_3253, n_3254, n_3255, 
      n_3256, n_3257, n_3258, n_3259, n_3260, n_3261, n_3262, n_3263, n_3264, 
      n_3265, n_3266, n_3267, n_3268, n_3269, n_3270, n_3271, n_3272, n_3273, 
      n_3274, n_3275, n_3276, n_3277, n_3278, n_3279, n_3280, n_3281, n_3282, 
      n_3283, n_3284, n_3285, n_3286, n_3287, n_3288, n_3289, n_3290, n_3291, 
      n_3292, n_3293, n_3294, n_3295, n_3296, n_3297, n_3298, n_3299, n_3300, 
      n_3301, n_3302, n_3303, n_3304, n_3305, n_3306, n_3307, n_3308, n_3309, 
      n_3310, n_3311, n_3312, n_3313, n_3314, n_3315, n_3316, n_3317, n_3318, 
      n_3319, n_3320, n_3321, n_3322, n_3323, n_3324, n_3325, n_3326, n_3327, 
      n_3328, n_3329, n_3330, n_3331, n_3332, n_3333, n_3334, n_3335, n_3336, 
      n_3337, n_3338, n_3339, n_3340, n_3341, n_3342, n_3343, n_3344, n_3345, 
      n_3346, n_3347, n_3348, n_3349, n_3350, n_3351, n_3352, n_3353, n_3354, 
      n_3355, n_3356, n_3357, n_3358, n_3359, n_3360, n_3361, n_3362, n_3363, 
      n_3364, n_3365, n_3366, n_3367, n_3368, n_3369, n_3370, n_3371, n_3372, 
      n_3373, n_3374, n_3375, n_3376, n_3377, n_3378, n_3379, n_3380, n_3381, 
      n_3382, n_3383, n_3384, n_3385, n_3386, n_3387, n_3388, n_3389, n_3390, 
      n_3391, n_3392, n_3393, n_3394, n_3395, n_3396, n_3397, n_3398, n_3399, 
      n_3400, n_3401, n_3402, n_3403, n_3404, n_3405, n_3406, n_3407, n_3408, 
      n_3409, n_3410, n_3411, n_3412, n_3413, n_3414, n_3415, n_3416, n_3417, 
      n_3418, n_3419, n_3420, n_3421, n_3422, n_3423, n_3424, n_3425 : 
      std_logic;

begin
   DATA_O <= ( DATA_O_7_port, DATA_O_6_port, DATA_O_5_port, DATA_O_4_port, 
      DATA_O_3_port, DATA_O_2_port, DATA_O_1_port, DATA_O_0_port );
   
   GET_KEY_reg : FD1 port map( D => N192, CP => CLK_I, Q => GET_KEY, QN => 
                           n3949);
   v_CNT4_reg_0_inst : FD1 port map( D => n4346, CP => CLK_I, Q => 
                           v_CNT4_0_port, QN => n4395);
   v_DATA_COLUMN_reg_24_inst : FD1 port map( D => n4837, CP => CLK_I, Q => 
                           v_DATA_COLUMN_24_port, QN => n_3156);
   v_DATA_COLUMN_reg_25_inst : FD1 port map( D => n4833, CP => CLK_I, Q => 
                           v_DATA_COLUMN_25_port, QN => n_3157);
   v_DATA_COLUMN_reg_26_inst : FD1 port map( D => n4829, CP => CLK_I, Q => 
                           v_DATA_COLUMN_26_port, QN => n_3158);
   v_DATA_COLUMN_reg_27_inst : FD1 port map( D => n4825, CP => CLK_I, Q => 
                           v_DATA_COLUMN_27_port, QN => n_3159);
   v_DATA_COLUMN_reg_28_inst : FD1 port map( D => n4821, CP => CLK_I, Q => 
                           v_DATA_COLUMN_28_port, QN => n_3160);
   v_DATA_COLUMN_reg_29_inst : FD1 port map( D => n4817, CP => CLK_I, Q => 
                           v_DATA_COLUMN_29_port, QN => n_3161);
   v_DATA_COLUMN_reg_30_inst : FD1 port map( D => n4813, CP => CLK_I, Q => 
                           v_DATA_COLUMN_30_port, QN => n_3162);
   v_DATA_COLUMN_reg_31_inst : FD1 port map( D => n4809, CP => CLK_I, Q => 
                           v_DATA_COLUMN_31_port, QN => n_3163);
   v_CNT4_reg_1_inst : FD1 port map( D => n4337, CP => CLK_I, Q => 
                           v_CNT4_1_port, QN => n4426);
   v_DATA_COLUMN_reg_8_inst : FD1 port map( D => n4836, CP => CLK_I, Q => 
                           v_DATA_COLUMN_8_port, QN => n_3164);
   v_DATA_COLUMN_reg_9_inst : FD1 port map( D => n4832, CP => CLK_I, Q => 
                           v_DATA_COLUMN_9_port, QN => n_3165);
   v_DATA_COLUMN_reg_10_inst : FD1 port map( D => n4831, CP => CLK_I, Q => 
                           v_DATA_COLUMN_10_port, QN => n_3166);
   v_DATA_COLUMN_reg_11_inst : FD1 port map( D => n4827, CP => CLK_I, Q => 
                           v_DATA_COLUMN_11_port, QN => n_3167);
   v_DATA_COLUMN_reg_12_inst : FD1 port map( D => n4823, CP => CLK_I, Q => 
                           v_DATA_COLUMN_12_port, QN => n_3168);
   v_DATA_COLUMN_reg_13_inst : FD1 port map( D => n4819, CP => CLK_I, Q => 
                           v_DATA_COLUMN_13_port, QN => n_3169);
   v_DATA_COLUMN_reg_14_inst : FD1 port map( D => n4815, CP => CLK_I, Q => 
                           v_DATA_COLUMN_14_port, QN => n_3170);
   v_DATA_COLUMN_reg_15_inst : FD1 port map( D => n4811, CP => CLK_I, Q => 
                           v_DATA_COLUMN_15_port, QN => n_3171);
   v_DATA_COLUMN_reg_16_inst : FD1 port map( D => n4838, CP => CLK_I, Q => 
                           v_DATA_COLUMN_16_port, QN => n_3172);
   v_DATA_COLUMN_reg_17_inst : FD1 port map( D => n4835, CP => CLK_I, Q => 
                           v_DATA_COLUMN_17_port, QN => n_3173);
   v_DATA_COLUMN_reg_18_inst : FD1 port map( D => n4830, CP => CLK_I, Q => 
                           v_DATA_COLUMN_18_port, QN => n_3174);
   v_DATA_COLUMN_reg_19_inst : FD1 port map( D => n4826, CP => CLK_I, Q => 
                           v_DATA_COLUMN_19_port, QN => n_3175);
   v_DATA_COLUMN_reg_20_inst : FD1 port map( D => n4822, CP => CLK_I, Q => 
                           v_DATA_COLUMN_20_port, QN => n_3176);
   v_DATA_COLUMN_reg_21_inst : FD1 port map( D => n4818, CP => CLK_I, Q => 
                           v_DATA_COLUMN_21_port, QN => n_3177);
   v_DATA_COLUMN_reg_22_inst : FD1 port map( D => n4814, CP => CLK_I, Q => 
                           v_DATA_COLUMN_22_port, QN => n_3178);
   v_DATA_COLUMN_reg_23_inst : FD1 port map( D => n4810, CP => CLK_I, Q => 
                           v_DATA_COLUMN_23_port, QN => n_3179);
   v_DATA_COLUMN_reg_0_inst : FD1 port map( D => n4839, CP => CLK_I, Q => 
                           v_DATA_COLUMN_0_port, QN => n_3180);
   v_DATA_COLUMN_reg_1_inst : FD1 port map( D => n4834, CP => CLK_I, Q => 
                           v_DATA_COLUMN_1_port, QN => n_3181);
   v_DATA_COLUMN_reg_2_inst : FD1 port map( D => n4828, CP => CLK_I, Q => 
                           v_DATA_COLUMN_2_port, QN => n_3182);
   v_DATA_COLUMN_reg_3_inst : FD1 port map( D => n4824, CP => CLK_I, Q => 
                           v_DATA_COLUMN_3_port, QN => n_3183);
   v_DATA_COLUMN_reg_4_inst : FD1 port map( D => n4820, CP => CLK_I, Q => 
                           v_DATA_COLUMN_4_port, QN => n_3184);
   v_DATA_COLUMN_reg_5_inst : FD1 port map( D => n4816, CP => CLK_I, Q => 
                           v_DATA_COLUMN_5_port, QN => n_3185);
   v_DATA_COLUMN_reg_6_inst : FD1 port map( D => n4812, CP => CLK_I, Q => 
                           v_DATA_COLUMN_6_port, QN => n_3186);
   v_DATA_COLUMN_reg_7_inst : FD1 port map( D => n4808, CP => CLK_I, Q => 
                           v_DATA_COLUMN_7_port, QN => n_3187);
   FF_VALID_DATA_reg : FD1 port map( D => n4312, CP => CLK_I, Q => n4527, QN =>
                           n3956);
   LAST_ROUND_reg : FD1 port map( D => n4311, CP => CLK_I, Q => n4441, QN => 
                           n3955);
   v_CALCULATION_CNTR_reg_0_inst : FD1 port map( D => n4310, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_0_port, QN => n4601);
   v_CALCULATION_CNTR_reg_1_inst : FD1 port map( D => n4309, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_1_port, QN => n4407);
   v_CALCULATION_CNTR_reg_2_inst : FD1 port map( D => n4308, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_2_port, QN => n4579);
   v_CALCULATION_CNTR_reg_3_inst : FD1 port map( D => n4307, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_3_port, QN => n4384);
   v_CALCULATION_CNTR_reg_4_inst : FD1 port map( D => n4306, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_4_port, QN => n4502);
   v_CALCULATION_CNTR_reg_5_inst : FD1 port map( D => n4848, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_5_port, QN => n_3188);
   v_CALCULATION_CNTR_reg_6_inst : FD1 port map( D => n4847, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_6_port, QN => n4600);
   v_CALCULATION_CNTR_reg_7_inst : FD1 port map( D => n4846, CP => CLK_I, Q => 
                           v_CALCULATION_CNTR_7_port, QN => n_3189);
   FF_GET_KEY_reg : FD1 port map( D => n4302, CP => CLK_I, Q => n_3190, QN => 
                           n3948);
   SRAM_WREN0_reg : FD1 port map( D => n4301, CP => CLK_I, Q => n_3191, QN => 
                           n3947);
   i_RAM_ADDR_WR0_reg_0_inst : FD1 port map( D => n4300, CP => CLK_I, Q => 
                           n_3192, QN => n3946);
   i_RAM_ADDR_WR0_reg_1_inst : FD1 port map( D => n4842, CP => CLK_I, Q => 
                           n4462, QN => n3945);
   v_KEY_NUMB_reg_5_inst : FD1 port map( D => n4298, CP => CLK_I, Q => 
                           v_INV_KEY_NUMB_5_port, QN => n3944);
   v_KEY_NUMB_reg_0_inst : FD1 port map( D => n4297, CP => CLK_I, Q => n_3193, 
                           QN => n4620);
   v_KEY_NUMB_reg_1_inst : FD1 port map( D => n4296, CP => CLK_I, Q => n_3194, 
                           QN => n4653);
   v_KEY_NUMB_reg_2_inst : FD1 port map( D => n4295, CP => CLK_I, Q => 
                           v_INV_KEY_NUMB_2_port, QN => n3943);
   v_KEY_NUMB_reg_3_inst : FD1 port map( D => n4294, CP => CLK_I, Q => 
                           v_INV_KEY_NUMB_3_port, QN => n3942);
   v_KEY_NUMB_reg_4_inst : FD1 port map( D => n4293, CP => CLK_I, Q => 
                           v_INV_KEY_NUMB_4_port, QN => n3941);
   i_RAM_ADDR_RD0_reg_0_inst : FD1 port map( D => n4292, CP => CLK_I, Q => 
                           n4602, QN => n3940);
   i_RAM_ADDR_RD0_reg_1_inst : FD1 port map( D => n4291, CP => CLK_I, Q => 
                           n4380, QN => n3939);
   CALCULATION_reg : FD1 port map( D => n4290, CP => CLK_I, Q => n_3195, QN => 
                           n3954);
   i_ROUND_reg_0_inst : FD1 port map( D => n4289, CP => CLK_I, Q => n_3196, QN 
                           => n3951);
   i_ROUND_reg_1_inst : FD1 port map( D => n4288, CP => CLK_I, Q => n4463, QN 
                           => n3950);
   i_ROUND_reg_2_inst : FD1 port map( D => n4287, CP => CLK_I, Q => n4619, QN 
                           => n3952);
   i_ROUND_reg_3_inst : FD1 port map( D => n4286, CP => CLK_I, Q => n_3197, QN 
                           => n3953);
   STATE_TABLE1_reg_0_7_inst : FD1 port map( D => n4285, CP => CLK_I, Q => 
                           n4417, QN => n_3198);
   STATE_TABLE1_reg_0_6_inst : FD1 port map( D => n4284, CP => CLK_I, Q => 
                           n4416, QN => n_3199);
   STATE_TABLE1_reg_0_5_inst : FD1 port map( D => n4283, CP => CLK_I, Q => 
                           n4604, QN => n3936);
   STATE_TABLE1_reg_0_4_inst : FD1 port map( D => n4282, CP => CLK_I, Q => 
                           n4547, QN => n_3200);
   STATE_TABLE1_reg_0_3_inst : FD1 port map( D => n4281, CP => CLK_I, Q => 
                           n4546, QN => n_3201);
   STATE_TABLE1_reg_0_2_inst : FD1 port map( D => n4280, CP => CLK_I, Q => 
                           n4517, QN => n_3202);
   STATE_TABLE1_reg_0_1_inst : FD1 port map( D => n4279, CP => CLK_I, Q => 
                           n4603, QN => n3932);
   STATE_TABLE1_reg_0_0_inst : FD1 port map( D => n4278, CP => CLK_I, Q => 
                           n4545, QN => n_3203);
   STATE_TABLE1_reg_1_7_inst : FD1 port map( D => n4277, CP => CLK_I, Q => 
                           n4607, QN => n3930);
   STATE_TABLE1_reg_1_6_inst : FD1 port map( D => n4276, CP => CLK_I, Q => 
                           n4431, QN => n_3204);
   STATE_TABLE1_reg_1_5_inst : FD1 port map( D => n4275, CP => CLK_I, Q => 
                           n4606, QN => n3928);
   STATE_TABLE1_reg_1_4_inst : FD1 port map( D => n4274, CP => CLK_I, Q => 
                           n4550, QN => n_3205);
   STATE_TABLE1_reg_1_3_inst : FD1 port map( D => n4273, CP => CLK_I, Q => 
                           n4444, QN => n_3206);
   STATE_TABLE1_reg_1_2_inst : FD1 port map( D => n4272, CP => CLK_I, Q => 
                           n4532, QN => n_3207);
   STATE_TABLE1_reg_1_1_inst : FD1 port map( D => n4271, CP => CLK_I, Q => 
                           n4605, QN => n3924);
   STATE_TABLE1_reg_1_0_inst : FD1 port map( D => n4270, CP => CLK_I, Q => 
                           n4519, QN => n_3208);
   STATE_TABLE1_reg_2_7_inst : FD1 port map( D => n4269, CP => CLK_I, Q => 
                           n4525, QN => n3922);
   STATE_TABLE1_reg_2_6_inst : FD1 port map( D => n4268, CP => CLK_I, Q => 
                           n4614, QN => n3921);
   STATE_TABLE1_reg_2_5_inst : FD1 port map( D => n4267, CP => CLK_I, Q => 
                           n4524, QN => n3920);
   STATE_TABLE1_reg_2_4_inst : FD1 port map( D => n4266, CP => CLK_I, Q => 
                           n4613, QN => n3919);
   STATE_TABLE1_reg_2_3_inst : FD1 port map( D => n4265, CP => CLK_I, Q => 
                           n4540, QN => n3918);
   STATE_TABLE1_reg_2_2_inst : FD1 port map( D => n4264, CP => CLK_I, Q => 
                           n4539, QN => n3917);
   STATE_TABLE1_reg_2_1_inst : FD1 port map( D => n4263, CP => CLK_I, Q => 
                           n4568, QN => n3916);
   STATE_TABLE1_reg_2_0_inst : FD1 port map( D => n4262, CP => CLK_I, Q => 
                           n4523, QN => n3915);
   STATE_TABLE1_reg_3_7_inst : FD1 port map( D => n4261, CP => CLK_I, Q => 
                           n4616, QN => n3914);
   STATE_TABLE1_reg_3_6_inst : FD1 port map( D => n4260, CP => CLK_I, Q => 
                           n4438, QN => n3913);
   STATE_TABLE1_reg_3_5_inst : FD1 port map( D => n4259, CP => CLK_I, Q => 
                           n4510, QN => n3912);
   STATE_TABLE1_reg_3_4_inst : FD1 port map( D => n4258, CP => CLK_I, Q => 
                           n4615, QN => n3911);
   STATE_TABLE1_reg_3_3_inst : FD1 port map( D => n4257, CP => CLK_I, Q => 
                           n4451, QN => n3910);
   STATE_TABLE1_reg_3_2_inst : FD1 port map( D => n4256, CP => CLK_I, Q => 
                           n4541, QN => n3909);
   STATE_TABLE1_reg_3_1_inst : FD1 port map( D => n4255, CP => CLK_I, Q => 
                           n4560, QN => n3908);
   STATE_TABLE1_reg_3_0_inst : FD1 port map( D => n4254, CP => CLK_I, Q => 
                           n4456, QN => n3907);
   STATE_TABLE1_reg_4_7_inst : FD1 port map( D => n4253, CP => CLK_I, Q => 
                           n4439, QN => n3906);
   STATE_TABLE1_reg_4_6_inst : FD1 port map( D => n4252, CP => CLK_I, Q => 
                           n4425, QN => n3905);
   STATE_TABLE1_reg_4_5_inst : FD1 port map( D => n4251, CP => CLK_I, Q => 
                           n4618, QN => n3904);
   STATE_TABLE1_reg_4_4_inst : FD1 port map( D => n4250, CP => CLK_I, Q => 
                           n4563, QN => n3903);
   STATE_TABLE1_reg_4_3_inst : FD1 port map( D => n4249, CP => CLK_I, Q => 
                           n4562, QN => n3902);
   STATE_TABLE1_reg_4_2_inst : FD1 port map( D => n4248, CP => CLK_I, Q => 
                           n4542, QN => n3901);
   STATE_TABLE1_reg_4_1_inst : FD1 port map( D => n4247, CP => CLK_I, Q => 
                           n4617, QN => n3900);
   STATE_TABLE1_reg_4_0_inst : FD1 port map( D => n4246, CP => CLK_I, Q => 
                           n4561, QN => n3899);
   STATE_TABLE1_reg_5_7_inst : FD1 port map( D => n4245, CP => CLK_I, Q => 
                           n4581, QN => n3898);
   STATE_TABLE1_reg_5_6_inst : FD1 port map( D => n4244, CP => CLK_I, Q => 
                           n4433, QN => n_3209);
   STATE_TABLE1_reg_5_5_inst : FD1 port map( D => n4243, CP => CLK_I, Q => 
                           n4580, QN => n3896);
   STATE_TABLE1_reg_5_4_inst : FD1 port map( D => n4242, CP => CLK_I, Q => 
                           n4446, QN => n_3210);
   STATE_TABLE1_reg_5_3_inst : FD1 port map( D => n4241, CP => CLK_I, Q => 
                           n4455, QN => n_3211);
   STATE_TABLE1_reg_5_2_inst : FD1 port map( D => n4240, CP => CLK_I, Q => 
                           n4432, QN => n_3212);
   STATE_TABLE1_reg_5_1_inst : FD1 port map( D => n4239, CP => CLK_I, Q => 
                           n4445, QN => n_3213);
   STATE_TABLE1_reg_5_0_inst : FD1 port map( D => n4238, CP => CLK_I, Q => 
                           n4419, QN => n_3214);
   STATE_TABLE1_reg_6_7_inst : FD1 port map( D => n4237, CP => CLK_I, Q => 
                           n4420, QN => n_3215);
   STATE_TABLE1_reg_6_6_inst : FD1 port map( D => n4236, CP => CLK_I, Q => 
                           n4583, QN => n3889);
   STATE_TABLE1_reg_6_5_inst : FD1 port map( D => n4235, CP => CLK_I, Q => 
                           n4415, QN => n_3216);
   STATE_TABLE1_reg_6_4_inst : FD1 port map( D => n4234, CP => CLK_I, Q => 
                           n4582, QN => n3887);
   STATE_TABLE1_reg_6_3_inst : FD1 port map( D => n4233, CP => CLK_I, Q => 
                           n4552, QN => n_3217);
   STATE_TABLE1_reg_6_2_inst : FD1 port map( D => n4232, CP => CLK_I, Q => 
                           n4551, QN => n_3218);
   STATE_TABLE1_reg_6_1_inst : FD1 port map( D => n4231, CP => CLK_I, Q => 
                           n4570, QN => n_3219);
   STATE_TABLE1_reg_6_0_inst : FD1 port map( D => n4230, CP => CLK_I, Q => 
                           n4520, QN => n_3220);
   STATE_TABLE1_reg_7_7_inst : FD1 port map( D => n4229, CP => CLK_I, Q => 
                           n4591, QN => n3882);
   STATE_TABLE1_reg_7_6_inst : FD1 port map( D => n4228, CP => CLK_I, Q => 
                           n4427, QN => n_3221);
   STATE_TABLE1_reg_7_5_inst : FD1 port map( D => n4227, CP => CLK_I, Q => 
                           n4507, QN => n_3222);
   STATE_TABLE1_reg_7_4_inst : FD1 port map( D => n4226, CP => CLK_I, Q => 
                           n4590, QN => n3879);
   STATE_TABLE1_reg_7_3_inst : FD1 port map( D => n4225, CP => CLK_I, Q => 
                           n4453, QN => n_3223);
   STATE_TABLE1_reg_7_2_inst : FD1 port map( D => n4224, CP => CLK_I, Q => 
                           n4544, QN => n_3224);
   STATE_TABLE1_reg_7_1_inst : FD1 port map( D => n4223, CP => CLK_I, Q => 
                           n4543, QN => n_3225);
   STATE_TABLE1_reg_7_0_inst : FD1 port map( D => n4222, CP => CLK_I, Q => 
                           n4440, QN => n_3226);
   STATE_TABLE1_reg_8_7_inst : FD1 port map( D => n4221, CP => CLK_I, Q => 
                           n4422, QN => n_3227);
   STATE_TABLE1_reg_8_6_inst : FD1 port map( D => n4220, CP => CLK_I, Q => 
                           n4397, QN => n_3228);
   STATE_TABLE1_reg_8_5_inst : FD1 port map( D => n4219, CP => CLK_I, Q => 
                           n4596, QN => n3872);
   STATE_TABLE1_reg_8_4_inst : FD1 port map( D => n4218, CP => CLK_I, Q => 
                           n4447, QN => n_3229);
   STATE_TABLE1_reg_8_3_inst : FD1 port map( D => n4217, CP => CLK_I, Q => 
                           n4554, QN => n_3230);
   STATE_TABLE1_reg_8_2_inst : FD1 port map( D => n4216, CP => CLK_I, Q => 
                           n4421, QN => n_3231);
   STATE_TABLE1_reg_8_1_inst : FD1 port map( D => n4215, CP => CLK_I, Q => 
                           n4595, QN => n3868);
   STATE_TABLE1_reg_8_0_inst : FD1 port map( D => n4214, CP => CLK_I, Q => 
                           n4553, QN => n_3232);
   STATE_TABLE1_reg_9_7_inst : FD1 port map( D => n4213, CP => CLK_I, Q => 
                           n4599, QN => n3866);
   STATE_TABLE1_reg_9_6_inst : FD1 port map( D => n4212, CP => CLK_I, Q => 
                           n4434, QN => n_3233);
   STATE_TABLE1_reg_9_5_inst : FD1 port map( D => n4211, CP => CLK_I, Q => 
                           n4598, QN => n3864);
   STATE_TABLE1_reg_9_4_inst : FD1 port map( D => n4210, CP => CLK_I, Q => 
                           n4449, QN => n_3234);
   STATE_TABLE1_reg_9_3_inst : FD1 port map( D => n4209, CP => CLK_I, Q => 
                           n4448, QN => n_3235);
   STATE_TABLE1_reg_9_2_inst : FD1 port map( D => n4208, CP => CLK_I, Q => 
                           n4533, QN => n_3236);
   STATE_TABLE1_reg_9_1_inst : FD1 port map( D => n4207, CP => CLK_I, Q => 
                           n4597, QN => n3860);
   STATE_TABLE1_reg_9_0_inst : FD1 port map( D => n4206, CP => CLK_I, Q => 
                           n4423, QN => n_3237);
   STATE_TABLE1_reg_10_7_inst : FD1 port map( D => n4205, CP => CLK_I, Q => 
                           n4522, QN => n3858);
   STATE_TABLE1_reg_10_6_inst : FD1 port map( D => n4204, CP => CLK_I, Q => 
                           n4609, QN => n3857);
   STATE_TABLE1_reg_10_5_inst : FD1 port map( D => n4203, CP => CLK_I, Q => 
                           n4521, QN => n3856);
   STATE_TABLE1_reg_10_4_inst : FD1 port map( D => n4202, CP => CLK_I, Q => 
                           n4608, QN => n3855);
   STATE_TABLE1_reg_10_3_inst : FD1 port map( D => n4201, CP => CLK_I, Q => 
                           n4536, QN => n3854);
   STATE_TABLE1_reg_10_2_inst : FD1 port map( D => n4200, CP => CLK_I, Q => 
                           n4535, QN => n3853);
   STATE_TABLE1_reg_10_1_inst : FD1 port map( D => n4199, CP => CLK_I, Q => 
                           n4567, QN => n3852);
   STATE_TABLE1_reg_10_0_inst : FD1 port map( D => n4198, CP => CLK_I, Q => 
                           n4534, QN => n3851);
   STATE_TABLE1_reg_11_7_inst : FD1 port map( D => n4197, CP => CLK_I, Q => 
                           n4593, QN => n3850);
   STATE_TABLE1_reg_11_6_inst : FD1 port map( D => n4196, CP => CLK_I, Q => 
                           n4428, QN => n_3238);
   STATE_TABLE1_reg_11_5_inst : FD1 port map( D => n4195, CP => CLK_I, Q => 
                           n4413, QN => n_3239);
   STATE_TABLE1_reg_11_4_inst : FD1 port map( D => n4194, CP => CLK_I, Q => 
                           n4592, QN => n3847);
   STATE_TABLE1_reg_11_3_inst : FD1 port map( D => n4193, CP => CLK_I, Q => 
                           n4443, QN => n_3240);
   STATE_TABLE1_reg_11_2_inst : FD1 port map( D => n4192, CP => CLK_I, Q => 
                           n4528, QN => n_3241);
   STATE_TABLE1_reg_11_1_inst : FD1 port map( D => n4191, CP => CLK_I, Q => 
                           n4442, QN => n_3242);
   STATE_TABLE1_reg_11_0_inst : FD1 port map( D => n4190, CP => CLK_I, Q => 
                           n4454, QN => n_3243);
   STATE_TABLE1_reg_12_7_inst : FD1 port map( D => n4189, CP => CLK_I, Q => 
                           n4435, QN => n3842);
   STATE_TABLE1_reg_12_6_inst : FD1 port map( D => n4188, CP => CLK_I, Q => 
                           n4424, QN => n3841);
   STATE_TABLE1_reg_12_5_inst : FD1 port map( D => n4187, CP => CLK_I, Q => 
                           n_3244, QN => n3840);
   STATE_TABLE1_reg_12_4_inst : FD1 port map( D => n4186, CP => CLK_I, Q => 
                           n4557, QN => n3839);
   STATE_TABLE1_reg_12_3_inst : FD1 port map( D => n4185, CP => CLK_I, Q => 
                           n4538, QN => n3838);
   STATE_TABLE1_reg_12_2_inst : FD1 port map( D => n4184, CP => CLK_I, Q => 
                           n4537, QN => n3837);
   STATE_TABLE1_reg_12_1_inst : FD1 port map( D => n4183, CP => CLK_I, Q => 
                           n4556, QN => n3836);
   STATE_TABLE1_reg_12_0_inst : FD1 port map( D => n4182, CP => CLK_I, Q => 
                           n4555, QN => n3835);
   STATE_TABLE1_reg_13_7_inst : FD1 port map( D => n4181, CP => CLK_I, Q => 
                           n4418, QN => n_3245);
   STATE_TABLE1_reg_13_6_inst : FD1 port map( D => n4180, CP => CLK_I, Q => 
                           n4398, QN => n_3246);
   STATE_TABLE1_reg_13_5_inst : FD1 port map( D => n4179, CP => CLK_I, Q => 
                           n4414, QN => n_3247);
   STATE_TABLE1_reg_13_4_inst : FD1 port map( D => n4178, CP => CLK_I, Q => 
                           n4566, QN => n_3248);
   STATE_TABLE1_reg_13_3_inst : FD1 port map( D => n4177, CP => CLK_I, Q => 
                           n4401, QN => n_3249);
   STATE_TABLE1_reg_13_2_inst : FD1 port map( D => n4176, CP => CLK_I, Q => 
                           n4430, QN => n_3250);
   STATE_TABLE1_reg_13_1_inst : FD1 port map( D => n4175, CP => CLK_I, Q => 
                           n4429, QN => n_3251);
   STATE_TABLE1_reg_13_0_inst : FD1 port map( D => n4174, CP => CLK_I, Q => 
                           n4529, QN => n_3252);
   STATE_TABLE1_reg_14_7_inst : FD1 port map( D => n4173, CP => CLK_I, Q => 
                           n4518, QN => n_3253);
   STATE_TABLE1_reg_14_6_inst : FD1 port map( D => n4172, CP => CLK_I, Q => 
                           n4526, QN => n3825);
   STATE_TABLE1_reg_14_5_inst : FD1 port map( D => n4171, CP => CLK_I, Q => 
                           n4514, QN => n3824);
   STATE_TABLE1_reg_14_4_inst : FD1 port map( D => n4170, CP => CLK_I, Q => 
                           n4594, QN => n3823);
   STATE_TABLE1_reg_14_3_inst : FD1 port map( D => n4169, CP => CLK_I, Q => 
                           n4531, QN => n_3254);
   STATE_TABLE1_reg_14_2_inst : FD1 port map( D => n4168, CP => CLK_I, Q => 
                           n4549, QN => n_3255);
   STATE_TABLE1_reg_14_1_inst : FD1 port map( D => n4167, CP => CLK_I, Q => 
                           n4548, QN => n_3256);
   STATE_TABLE1_reg_14_0_inst : FD1 port map( D => n4166, CP => CLK_I, Q => 
                           n4530, QN => n_3257);
   STATE_TABLE1_reg_15_7_inst : FD1 port map( D => n4165, CP => CLK_I, Q => 
                           n4612, QN => n3818);
   STATE_TABLE1_reg_15_6_inst : FD1 port map( D => n4164, CP => CLK_I, Q => 
                           n4437, QN => n3817);
   STATE_TABLE1_reg_15_5_inst : FD1 port map( D => n4163, CP => CLK_I, Q => 
                           n4611, QN => n3816);
   v_RAM_IN0_reg_24_inst : FD1 port map( D => n4162, CP => CLK_I, Q => n_3258, 
                           QN => n4495);
   t_STATE_RAM0_reg_0_24_inst : FD1 port map( D => n4161, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_24_port, QN => n_3259);
   t_STATE_RAM0_reg_1_24_inst : FD1 port map( D => n4160, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_24_port, QN => n_3260);
   t_STATE_RAM0_reg_2_24_inst : FD1 port map( D => n4159, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_24_port, QN => n_3261);
   t_STATE_RAM0_reg_3_24_inst : FD1 port map( D => n4158, CP => CLK_I, Q => 
                           n_3262, QN => n4652);
   v_RAM_OUT0_reg_24_inst : FD1 port map( D => n4157, CP => CLK_I, Q => 
                           v_RAM_OUT0_24_port, QN => n4394);
   STATE_TABLE1_reg_15_4_inst : FD1 port map( D => n4156, CP => CLK_I, Q => 
                           n4610, QN => n3815);
   v_RAM_IN0_reg_31_inst : FD1 port map( D => n4155, CP => CLK_I, Q => n_3263, 
                           QN => n4494);
   t_STATE_RAM0_reg_0_31_inst : FD1 port map( D => n4154, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_31_port, QN => n_3264);
   t_STATE_RAM0_reg_1_31_inst : FD1 port map( D => n4153, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_31_port, QN => n_3265);
   t_STATE_RAM0_reg_2_31_inst : FD1 port map( D => n4152, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_31_port, QN => n_3266);
   t_STATE_RAM0_reg_3_31_inst : FD1 port map( D => n4151, CP => CLK_I, Q => 
                           n_3267, QN => n4651);
   v_RAM_OUT0_reg_31_inst : FD1 port map( D => n4150, CP => CLK_I, Q => 
                           v_RAM_OUT0_31_port, QN => n4587);
   v_RAM_IN0_reg_23_inst : FD1 port map( D => n4149, CP => CLK_I, Q => n_3268, 
                           QN => n4493);
   t_STATE_RAM0_reg_0_23_inst : FD1 port map( D => n4148, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_23_port, QN => n_3269);
   t_STATE_RAM0_reg_1_23_inst : FD1 port map( D => n4147, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_23_port, QN => n_3270);
   t_STATE_RAM0_reg_2_23_inst : FD1 port map( D => n4146, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_23_port, QN => n_3271);
   t_STATE_RAM0_reg_3_23_inst : FD1 port map( D => n4145, CP => CLK_I, Q => 
                           n_3272, QN => n4650);
   v_RAM_OUT0_reg_23_inst : FD1 port map( D => n4144, CP => CLK_I, Q => 
                           v_RAM_OUT0_23_port, QN => n4578);
   v_RAM_IN0_reg_15_inst : FD1 port map( D => n4143, CP => CLK_I, Q => n_3273, 
                           QN => n4492);
   t_STATE_RAM0_reg_0_15_inst : FD1 port map( D => n4142, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_15_port, QN => n_3274);
   t_STATE_RAM0_reg_1_15_inst : FD1 port map( D => n4141, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_15_port, QN => n_3275);
   t_STATE_RAM0_reg_2_15_inst : FD1 port map( D => n4140, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_15_port, QN => n_3276);
   t_STATE_RAM0_reg_3_15_inst : FD1 port map( D => n4139, CP => CLK_I, Q => 
                           n_3277, QN => n4649);
   v_RAM_OUT0_reg_15_inst : FD1 port map( D => n4138, CP => CLK_I, Q => 
                           v_RAM_OUT0_15_port, QN => n4396);
   v_RAM_IN0_reg_7_inst : FD1 port map( D => n4137, CP => CLK_I, Q => n_3278, 
                           QN => n4491);
   t_STATE_RAM0_reg_0_7_inst : FD1 port map( D => n4136, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_7_port, QN => n_3279);
   t_STATE_RAM0_reg_1_7_inst : FD1 port map( D => n4135, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_7_port, QN => n_3280);
   t_STATE_RAM0_reg_2_7_inst : FD1 port map( D => n4134, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_7_port, QN => n_3281);
   t_STATE_RAM0_reg_3_7_inst : FD1 port map( D => n4133, CP => CLK_I, Q => 
                           n_3282, QN => n4648);
   v_RAM_OUT0_reg_7_inst : FD1 port map( D => n4132, CP => CLK_I, Q => 
                           v_RAM_OUT0_7_port, QN => n4588);
   STATE_TABLE1_reg_15_3_inst : FD1 port map( D => n4131, CP => CLK_I, Q => 
                           n4436, QN => n3814);
   v_RAM_IN0_reg_30_inst : FD1 port map( D => n4130, CP => CLK_I, Q => n_3283, 
                           QN => n4490);
   t_STATE_RAM0_reg_0_30_inst : FD1 port map( D => n4129, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_30_port, QN => n_3284);
   t_STATE_RAM0_reg_1_30_inst : FD1 port map( D => n4128, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_30_port, QN => n_3285);
   t_STATE_RAM0_reg_2_30_inst : FD1 port map( D => n4127, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_30_port, QN => n_3286);
   t_STATE_RAM0_reg_3_30_inst : FD1 port map( D => n4126, CP => CLK_I, Q => 
                           n_3287, QN => n4647);
   v_RAM_OUT0_reg_30_inst : FD1 port map( D => n4125, CP => CLK_I, Q => 
                           v_RAM_OUT0_30_port, QN => n4508);
   v_RAM_IN0_reg_22_inst : FD1 port map( D => n4124, CP => CLK_I, Q => n_3288, 
                           QN => n4489);
   t_STATE_RAM0_reg_0_22_inst : FD1 port map( D => n4123, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_22_port, QN => n_3289);
   t_STATE_RAM0_reg_1_22_inst : FD1 port map( D => n4122, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_22_port, QN => n_3290);
   t_STATE_RAM0_reg_2_22_inst : FD1 port map( D => n4121, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_22_port, QN => n_3291);
   t_STATE_RAM0_reg_3_22_inst : FD1 port map( D => n4120, CP => CLK_I, Q => 
                           n_3292, QN => n4646);
   v_RAM_OUT0_reg_22_inst : FD1 port map( D => n4119, CP => CLK_I, Q => 
                           v_RAM_OUT0_22_port, QN => n4501);
   v_RAM_IN0_reg_14_inst : FD1 port map( D => n4118, CP => CLK_I, Q => n_3293, 
                           QN => n4488);
   t_STATE_RAM0_reg_0_14_inst : FD1 port map( D => n4117, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_14_port, QN => n_3294);
   t_STATE_RAM0_reg_1_14_inst : FD1 port map( D => n4116, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_14_port, QN => n_3295);
   t_STATE_RAM0_reg_2_14_inst : FD1 port map( D => n4115, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_14_port, QN => n_3296);
   t_STATE_RAM0_reg_3_14_inst : FD1 port map( D => n4114, CP => CLK_I, Q => 
                           n_3297, QN => n4645);
   v_RAM_OUT0_reg_14_inst : FD1 port map( D => n4113, CP => CLK_I, Q => 
                           v_RAM_OUT0_14_port, QN => n4509);
   v_RAM_IN0_reg_6_inst : FD1 port map( D => n4112, CP => CLK_I, Q => n_3298, 
                           QN => n4487);
   t_STATE_RAM0_reg_0_6_inst : FD1 port map( D => n4111, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_6_port, QN => n_3299);
   t_STATE_RAM0_reg_1_6_inst : FD1 port map( D => n4110, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_6_port, QN => n_3300);
   t_STATE_RAM0_reg_2_6_inst : FD1 port map( D => n4109, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_6_port, QN => n_3301);
   t_STATE_RAM0_reg_3_6_inst : FD1 port map( D => n4108, CP => CLK_I, Q => 
                           n_3302, QN => n4644);
   v_RAM_OUT0_reg_6_inst : FD1 port map( D => n4107, CP => CLK_I, Q => 
                           v_RAM_OUT0_6_port, QN => n4500);
   STATE_TABLE1_reg_15_2_inst : FD1 port map( D => n4106, CP => CLK_I, Q => 
                           n4559, QN => n3813);
   v_RAM_IN0_reg_21_inst : FD1 port map( D => n4105, CP => CLK_I, Q => n_3303, 
                           QN => n4486);
   t_STATE_RAM0_reg_0_21_inst : FD1 port map( D => n4104, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_21_port, QN => n_3304);
   t_STATE_RAM0_reg_1_21_inst : FD1 port map( D => n4103, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_21_port, QN => n_3305);
   t_STATE_RAM0_reg_2_21_inst : FD1 port map( D => n4102, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_21_port, QN => n_3306);
   t_STATE_RAM0_reg_3_21_inst : FD1 port map( D => n4101, CP => CLK_I, Q => 
                           n_3307, QN => n4643);
   v_RAM_OUT0_reg_21_inst : FD1 port map( D => n4100, CP => CLK_I, Q => 
                           v_RAM_OUT0_21_port, QN => n4409);
   v_RAM_IN0_reg_13_inst : FD1 port map( D => n4099, CP => CLK_I, Q => n_3308, 
                           QN => n4485);
   t_STATE_RAM0_reg_0_13_inst : FD1 port map( D => n4098, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_13_port, QN => n_3309);
   t_STATE_RAM0_reg_1_13_inst : FD1 port map( D => n4097, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_13_port, QN => n_3310);
   t_STATE_RAM0_reg_2_13_inst : FD1 port map( D => n4096, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_13_port, QN => n_3311);
   t_STATE_RAM0_reg_3_13_inst : FD1 port map( D => n4095, CP => CLK_I, Q => 
                           n_3312, QN => n4642);
   v_RAM_OUT0_reg_13_inst : FD1 port map( D => n4094, CP => CLK_I, Q => 
                           v_RAM_OUT0_13_port, QN => n4516);
   v_RAM_IN0_reg_29_inst : FD1 port map( D => n4093, CP => CLK_I, Q => n_3313, 
                           QN => n4484);
   t_STATE_RAM0_reg_0_29_inst : FD1 port map( D => n4092, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_29_port, QN => n_3314);
   t_STATE_RAM0_reg_1_29_inst : FD1 port map( D => n4091, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_29_port, QN => n_3315);
   t_STATE_RAM0_reg_2_29_inst : FD1 port map( D => n4090, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_29_port, QN => n_3316);
   t_STATE_RAM0_reg_3_29_inst : FD1 port map( D => n4089, CP => CLK_I, Q => 
                           n_3317, QN => n4641);
   v_RAM_OUT0_reg_29_inst : FD1 port map( D => n4088, CP => CLK_I, Q => 
                           v_RAM_OUT0_29_port, QN => n4410);
   v_RAM_IN0_reg_5_inst : FD1 port map( D => n4087, CP => CLK_I, Q => n_3318, 
                           QN => n4483);
   t_STATE_RAM0_reg_0_5_inst : FD1 port map( D => n4086, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_5_port, QN => n_3319);
   t_STATE_RAM0_reg_1_5_inst : FD1 port map( D => n4085, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_5_port, QN => n_3320);
   t_STATE_RAM0_reg_2_5_inst : FD1 port map( D => n4084, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_5_port, QN => n_3321);
   t_STATE_RAM0_reg_3_5_inst : FD1 port map( D => n4083, CP => CLK_I, Q => 
                           n_3322, QN => n4640);
   v_RAM_OUT0_reg_5_inst : FD1 port map( D => n4082, CP => CLK_I, Q => 
                           v_RAM_OUT0_5_port, QN => n4408);
   v_RAM_IN0_reg_2_inst : FD1 port map( D => n4081, CP => CLK_I, Q => n_3323, 
                           QN => n4482);
   t_STATE_RAM0_reg_0_2_inst : FD1 port map( D => n4080, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_2_port, QN => n_3324);
   t_STATE_RAM0_reg_1_2_inst : FD1 port map( D => n4079, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_2_port, QN => n_3325);
   t_STATE_RAM0_reg_2_2_inst : FD1 port map( D => n4078, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_2_port, QN => n_3326);
   t_STATE_RAM0_reg_3_2_inst : FD1 port map( D => n4077, CP => CLK_I, Q => 
                           n_3327, QN => n4639);
   v_RAM_OUT0_reg_2_inst : FD1 port map( D => n4076, CP => CLK_I, Q => 
                           v_RAM_OUT0_2_port, QN => n4363);
   STATE_TABLE1_reg_15_1_inst : FD1 port map( D => n4075, CP => CLK_I, Q => 
                           n4558, QN => n3812);
   v_RAM_IN0_reg_18_inst : FD1 port map( D => n4074, CP => CLK_I, Q => n_3328, 
                           QN => n4481);
   t_STATE_RAM0_reg_0_18_inst : FD1 port map( D => n4073, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_18_port, QN => n_3329);
   t_STATE_RAM0_reg_1_18_inst : FD1 port map( D => n4072, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_18_port, QN => n_3330);
   t_STATE_RAM0_reg_2_18_inst : FD1 port map( D => n4071, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_18_port, QN => n_3331);
   t_STATE_RAM0_reg_3_18_inst : FD1 port map( D => n4070, CP => CLK_I, Q => 
                           n_3332, QN => n4638);
   v_RAM_OUT0_reg_18_inst : FD1 port map( D => n4069, CP => CLK_I, Q => 
                           v_RAM_OUT0_18_port, QN => n4365);
   v_RAM_IN0_reg_28_inst : FD1 port map( D => n4068, CP => CLK_I, Q => n_3333, 
                           QN => n4480);
   t_STATE_RAM0_reg_0_28_inst : FD1 port map( D => n4067, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_28_port, QN => n_3334);
   t_STATE_RAM0_reg_1_28_inst : FD1 port map( D => n4066, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_28_port, QN => n_3335);
   t_STATE_RAM0_reg_2_28_inst : FD1 port map( D => n4065, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_28_port, QN => n_3336);
   t_STATE_RAM0_reg_3_28_inst : FD1 port map( D => n4064, CP => CLK_I, Q => 
                           n_3337, QN => n4637);
   v_RAM_OUT0_reg_28_inst : FD1 port map( D => n4063, CP => CLK_I, Q => 
                           v_RAM_OUT0_28_port, QN => n4368);
   v_RAM_IN0_reg_12_inst : FD1 port map( D => n4062, CP => CLK_I, Q => n_3338, 
                           QN => n4479);
   t_STATE_RAM0_reg_0_12_inst : FD1 port map( D => n4061, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_12_port, QN => n_3339);
   t_STATE_RAM0_reg_1_12_inst : FD1 port map( D => n4060, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_12_port, QN => n_3340);
   t_STATE_RAM0_reg_2_12_inst : FD1 port map( D => n4059, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_12_port, QN => n_3341);
   t_STATE_RAM0_reg_3_12_inst : FD1 port map( D => n4058, CP => CLK_I, Q => 
                           n_3342, QN => n4636);
   v_RAM_OUT0_reg_12_inst : FD1 port map( D => n4057, CP => CLK_I, Q => 
                           v_RAM_OUT0_12_port, QN => n4404);
   v_RAM_IN0_reg_20_inst : FD1 port map( D => n4056, CP => CLK_I, Q => n_3343, 
                           QN => n4478);
   t_STATE_RAM0_reg_0_20_inst : FD1 port map( D => n4055, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_20_port, QN => n_3344);
   t_STATE_RAM0_reg_1_20_inst : FD1 port map( D => n4054, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_20_port, QN => n_3345);
   t_STATE_RAM0_reg_2_20_inst : FD1 port map( D => n4053, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_20_port, QN => n_3346);
   t_STATE_RAM0_reg_3_20_inst : FD1 port map( D => n4052, CP => CLK_I, Q => 
                           n_3347, QN => n4635);
   v_RAM_OUT0_reg_20_inst : FD1 port map( D => n4051, CP => CLK_I, Q => 
                           v_RAM_OUT0_20_port, QN => n4364);
   v_RAM_IN0_reg_4_inst : FD1 port map( D => n4050, CP => CLK_I, Q => n_3348, 
                           QN => n4477);
   t_STATE_RAM0_reg_0_4_inst : FD1 port map( D => n4049, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_4_port, QN => n_3349);
   t_STATE_RAM0_reg_1_4_inst : FD1 port map( D => n4048, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_4_port, QN => n_3350);
   t_STATE_RAM0_reg_2_4_inst : FD1 port map( D => n4047, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_4_port, QN => n_3351);
   t_STATE_RAM0_reg_3_4_inst : FD1 port map( D => n4046, CP => CLK_I, Q => 
                           n_3352, QN => n4634);
   v_RAM_OUT0_reg_4_inst : FD1 port map( D => n4045, CP => CLK_I, Q => 
                           v_RAM_OUT0_4_port, QN => n4367);
   v_RAM_IN0_reg_1_inst : FD1 port map( D => n4044, CP => CLK_I, Q => n_3353, 
                           QN => n4476);
   t_STATE_RAM0_reg_0_1_inst : FD1 port map( D => n4043, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_1_port, QN => n_3354);
   t_STATE_RAM0_reg_1_1_inst : FD1 port map( D => n4042, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_1_port, QN => n_3355);
   t_STATE_RAM0_reg_2_1_inst : FD1 port map( D => n4041, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_1_port, QN => n_3356);
   t_STATE_RAM0_reg_3_1_inst : FD1 port map( D => n4040, CP => CLK_I, Q => 
                           n_3357, QN => n4633);
   v_RAM_OUT0_reg_1_inst : FD1 port map( D => n4039, CP => CLK_I, Q => 
                           v_RAM_OUT0_1_port, QN => n4497);
   v_RAM_IN0_reg_9_inst : FD1 port map( D => n4038, CP => CLK_I, Q => n_3358, 
                           QN => n4475);
   t_STATE_RAM0_reg_0_9_inst : FD1 port map( D => n4037, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_9_port, QN => n_3359);
   t_STATE_RAM0_reg_1_9_inst : FD1 port map( D => n4036, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_9_port, QN => n_3360);
   t_STATE_RAM0_reg_2_9_inst : FD1 port map( D => n4035, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_9_port, QN => n_3361);
   t_STATE_RAM0_reg_3_9_inst : FD1 port map( D => n4034, CP => CLK_I, Q => 
                           n_3362, QN => n4632);
   v_RAM_OUT0_reg_9_inst : FD1 port map( D => n4033, CP => CLK_I, Q => 
                           v_RAM_OUT0_9_port, QN => n4569);
   STATE_TABLE1_reg_15_0_inst : FD1 port map( D => n4032, CP => CLK_I, Q => 
                           n4450, QN => n3811);
   v_RAM_IN0_reg_26_inst : FD1 port map( D => n4031, CP => CLK_I, Q => n_3363, 
                           QN => n4474);
   t_STATE_RAM0_reg_0_26_inst : FD1 port map( D => n4030, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_26_port, QN => n_3364);
   t_STATE_RAM0_reg_1_26_inst : FD1 port map( D => n4029, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_26_port, QN => n_3365);
   t_STATE_RAM0_reg_2_26_inst : FD1 port map( D => n4028, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_26_port, QN => n_3366);
   t_STATE_RAM0_reg_3_26_inst : FD1 port map( D => n4027, CP => CLK_I, Q => 
                           n_3367, QN => n4631);
   v_RAM_OUT0_reg_26_inst : FD1 port map( D => n4026, CP => CLK_I, Q => 
                           v_RAM_OUT0_26_port, QN => n4362);
   v_RAM_IN0_reg_10_inst : FD1 port map( D => n4025, CP => CLK_I, Q => n_3368, 
                           QN => n4473);
   t_STATE_RAM0_reg_0_10_inst : FD1 port map( D => n4024, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_10_port, QN => n_3369);
   t_STATE_RAM0_reg_1_10_inst : FD1 port map( D => n4023, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_10_port, QN => n_3370);
   t_STATE_RAM0_reg_2_10_inst : FD1 port map( D => n4022, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_10_port, QN => n_3371);
   t_STATE_RAM0_reg_3_10_inst : FD1 port map( D => n4021, CP => CLK_I, Q => 
                           n_3372, QN => n4630);
   v_RAM_OUT0_reg_10_inst : FD1 port map( D => n4020, CP => CLK_I, Q => 
                           v_RAM_OUT0_10_port, QN => n4378);
   v_RAM_IN0_reg_27_inst : FD1 port map( D => n4019, CP => CLK_I, Q => n_3373, 
                           QN => n4472);
   t_STATE_RAM0_reg_0_27_inst : FD1 port map( D => n4018, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_27_port, QN => n_3374);
   t_STATE_RAM0_reg_1_27_inst : FD1 port map( D => n4017, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_27_port, QN => n_3375);
   t_STATE_RAM0_reg_2_27_inst : FD1 port map( D => n4016, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_27_port, QN => n_3376);
   t_STATE_RAM0_reg_3_27_inst : FD1 port map( D => n4015, CP => CLK_I, Q => 
                           n_3377, QN => n4629);
   v_RAM_OUT0_reg_27_inst : FD1 port map( D => n4014, CP => CLK_I, Q => 
                           v_RAM_OUT0_27_port, QN => n4411);
   v_RAM_IN0_reg_19_inst : FD1 port map( D => n4013, CP => CLK_I, Q => n_3378, 
                           QN => n4471);
   t_STATE_RAM0_reg_0_19_inst : FD1 port map( D => n4012, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_19_port, QN => n_3379);
   t_STATE_RAM0_reg_1_19_inst : FD1 port map( D => n4011, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_19_port, QN => n_3380);
   t_STATE_RAM0_reg_2_19_inst : FD1 port map( D => n4010, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_19_port, QN => n_3381);
   t_STATE_RAM0_reg_3_19_inst : FD1 port map( D => n4009, CP => CLK_I, Q => 
                           n_3382, QN => n4628);
   v_RAM_OUT0_reg_19_inst : FD1 port map( D => n4008, CP => CLK_I, Q => 
                           v_RAM_OUT0_19_port, QN => n4406);
   v_RAM_IN0_reg_11_inst : FD1 port map( D => n4007, CP => CLK_I, Q => n_3383, 
                           QN => n4470);
   t_STATE_RAM0_reg_0_11_inst : FD1 port map( D => n4006, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_11_port, QN => n_3384);
   t_STATE_RAM0_reg_1_11_inst : FD1 port map( D => n4005, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_11_port, QN => n_3385);
   t_STATE_RAM0_reg_2_11_inst : FD1 port map( D => n4004, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_11_port, QN => n_3386);
   t_STATE_RAM0_reg_3_11_inst : FD1 port map( D => n4003, CP => CLK_I, Q => 
                           n_3387, QN => n4627);
   v_RAM_OUT0_reg_11_inst : FD1 port map( D => n4002, CP => CLK_I, Q => 
                           v_RAM_OUT0_11_port, QN => n4412);
   v_RAM_IN0_reg_3_inst : FD1 port map( D => n4001, CP => CLK_I, Q => n_3388, 
                           QN => n4469);
   t_STATE_RAM0_reg_0_3_inst : FD1 port map( D => n4000, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_3_port, QN => n_3389);
   t_STATE_RAM0_reg_1_3_inst : FD1 port map( D => n3999, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_3_port, QN => n_3390);
   t_STATE_RAM0_reg_2_3_inst : FD1 port map( D => n3998, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_3_port, QN => n_3391);
   t_STATE_RAM0_reg_3_3_inst : FD1 port map( D => n3997, CP => CLK_I, Q => 
                           n_3392, QN => n4626);
   v_RAM_OUT0_reg_3_inst : FD1 port map( D => n3996, CP => CLK_I, Q => 
                           v_RAM_OUT0_3_port, QN => n4405);
   v_RAM_IN0_reg_25_inst : FD1 port map( D => n3995, CP => CLK_I, Q => n_3393, 
                           QN => n4468);
   t_STATE_RAM0_reg_0_25_inst : FD1 port map( D => n3994, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_25_port, QN => n_3394);
   t_STATE_RAM0_reg_1_25_inst : FD1 port map( D => n3993, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_25_port, QN => n_3395);
   t_STATE_RAM0_reg_2_25_inst : FD1 port map( D => n3992, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_25_port, QN => n_3396);
   t_STATE_RAM0_reg_3_25_inst : FD1 port map( D => n3991, CP => CLK_I, Q => 
                           n_3397, QN => n4625);
   v_RAM_OUT0_reg_25_inst : FD1 port map( D => n3990, CP => CLK_I, Q => 
                           v_RAM_OUT0_25_port, QN => n4499);
   v_RAM_IN0_reg_17_inst : FD1 port map( D => n3989, CP => CLK_I, Q => n_3398, 
                           QN => n4467);
   t_STATE_RAM0_reg_0_17_inst : FD1 port map( D => n3988, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_17_port, QN => n_3399);
   t_STATE_RAM0_reg_1_17_inst : FD1 port map( D => n3987, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_17_port, QN => n_3400);
   t_STATE_RAM0_reg_2_17_inst : FD1 port map( D => n3986, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_17_port, QN => n_3401);
   t_STATE_RAM0_reg_3_17_inst : FD1 port map( D => n3985, CP => CLK_I, Q => 
                           n_3402, QN => n4624);
   v_RAM_OUT0_reg_17_inst : FD1 port map( D => n3984, CP => CLK_I, Q => 
                           v_RAM_OUT0_17_port, QN => n4498);
   v_RAM_IN0_reg_8_inst : FD1 port map( D => n3983, CP => CLK_I, Q => n_3403, 
                           QN => n4466);
   t_STATE_RAM0_reg_0_8_inst : FD1 port map( D => n3982, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_8_port, QN => n_3404);
   t_STATE_RAM0_reg_1_8_inst : FD1 port map( D => n3981, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_8_port, QN => n_3405);
   t_STATE_RAM0_reg_2_8_inst : FD1 port map( D => n3980, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_8_port, QN => n_3406);
   t_STATE_RAM0_reg_3_8_inst : FD1 port map( D => n3979, CP => CLK_I, Q => 
                           n_3407, QN => n4623);
   v_RAM_OUT0_reg_8_inst : FD1 port map( D => n3978, CP => CLK_I, Q => 
                           v_RAM_OUT0_8_port, QN => n4391);
   v_RAM_IN0_reg_16_inst : FD1 port map( D => n3977, CP => CLK_I, Q => n_3408, 
                           QN => n4465);
   t_STATE_RAM0_reg_0_16_inst : FD1 port map( D => n3976, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_16_port, QN => n_3409);
   t_STATE_RAM0_reg_1_16_inst : FD1 port map( D => n3975, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_16_port, QN => n_3410);
   t_STATE_RAM0_reg_2_16_inst : FD1 port map( D => n3974, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_16_port, QN => n_3411);
   t_STATE_RAM0_reg_3_16_inst : FD1 port map( D => n3973, CP => CLK_I, Q => 
                           n_3412, QN => n4622);
   v_RAM_OUT0_reg_16_inst : FD1 port map( D => n3972, CP => CLK_I, Q => 
                           v_RAM_OUT0_16_port, QN => n4393);
   v_RAM_IN0_reg_0_inst : FD1 port map( D => n3971, CP => CLK_I, Q => n_3413, 
                           QN => n4464);
   t_STATE_RAM0_reg_0_0_inst : FD1 port map( D => n3970, CP => CLK_I, Q => 
                           t_STATE_RAM0_0_0_port, QN => n_3414);
   t_STATE_RAM0_reg_1_0_inst : FD1 port map( D => n3969, CP => CLK_I, Q => 
                           t_STATE_RAM0_1_0_port, QN => n_3415);
   t_STATE_RAM0_reg_2_0_inst : FD1 port map( D => n3968, CP => CLK_I, Q => 
                           t_STATE_RAM0_2_0_port, QN => n_3416);
   t_STATE_RAM0_reg_3_0_inst : FD1 port map( D => n3967, CP => CLK_I, Q => 
                           n_3417, QN => n4621);
   v_RAM_OUT0_reg_0_inst : FD1 port map( D => n3966, CP => CLK_I, Q => 
                           v_RAM_OUT0_0_port, QN => n4392);
   DATA_O_reg_7_inst : FD1 port map( D => n3965, CP => CLK_I, Q => 
                           DATA_O_7_port, QN => n_3418);
   DATA_O_reg_6_inst : FD1 port map( D => n3964, CP => CLK_I, Q => 
                           DATA_O_6_port, QN => n_3419);
   DATA_O_reg_5_inst : FD1 port map( D => n3963, CP => CLK_I, Q => 
                           DATA_O_5_port, QN => n_3420);
   DATA_O_reg_4_inst : FD1 port map( D => n3962, CP => CLK_I, Q => 
                           DATA_O_4_port, QN => n_3421);
   DATA_O_reg_3_inst : FD1 port map( D => n3961, CP => CLK_I, Q => 
                           DATA_O_3_port, QN => n_3422);
   DATA_O_reg_2_inst : FD1 port map( D => n3960, CP => CLK_I, Q => 
                           DATA_O_2_port, QN => n_3423);
   DATA_O_reg_1_inst : FD1 port map( D => n3959, CP => CLK_I, Q => 
                           DATA_O_1_port, QN => n_3424);
   DATA_O_reg_0_inst : FD1 port map( D => n3958, CP => CLK_I, Q => 
                           DATA_O_0_port, QN => n_3425);
   VALID_O_reg : FD1 port map( D => n3957, CP => CLK_I, Q => VALID_O, QN => 
                           n3810);
   U1258 : AN3 port map( A => n4426, B => n4395, C => n4527, Z => n1353);
   U1259 : OR3 port map( A => n1351, B => n4860, C => n1391, Z => n1387);
   U1605 : AN3 port map( A => n1502, B => n1503, C => n1504, Z => n1501);
   U1615 : OR3 port map( A => n4388, B => n4599, C => n1527, Z => n1525);
   U1619 : OR3 port map( A => n4577, B => n4434, C => n1527, Z => n1532);
   U1623 : OR3 port map( A => n4385, B => n4598, C => n1527, Z => n1537);
   U1627 : OR3 port map( A => n4799, B => n4449, C => n1527, Z => n1542);
   U1631 : OR3 port map( A => n4576, B => n4448, C => n1527, Z => n1546);
   U1635 : OR3 port map( A => n4390, B => n4533, C => n1527, Z => n1551);
   U1639 : OR3 port map( A => n4725, B => n4597, C => n1527, Z => n1555);
   U1643 : OR3 port map( A => n4732, B => n4423, C => n1527, Z => n1560);
   U1649 : OR3 port map( A => n4575, B => n4422, C => n1527, Z => n1566);
   U1653 : OR3 port map( A => n4574, B => n4397, C => n1527, Z => n1572);
   U1657 : OR3 port map( A => n4461, B => n4596, C => n1527, Z => n1577);
   U1661 : OR3 port map( A => n4760, B => n4447, C => n1527, Z => n1583);
   U1665 : OR3 port map( A => n4761, B => n4554, C => n1527, Z => n1587);
   U1669 : OR3 port map( A => n4771, B => n4421, C => n1527, Z => n1591);
   U1673 : OR3 port map( A => n4787, B => n4595, C => n1527, Z => n1595);
   U1677 : OR3 port map( A => n4804, B => n4553, C => n1527, Z => n1600);
   U1683 : OR3 port map( A => n4459, B => n4591, C => n1609, Z => n1606);
   U1687 : OR3 port map( A => n4573, B => n4427, C => n1609, Z => n1614);
   U1691 : OR3 port map( A => n4773, B => n4507, C => n1609, Z => n1619);
   U1695 : OR3 port map( A => n4458, B => n4590, C => n1609, Z => n1623);
   U1699 : OR3 port map( A => n4572, B => n4453, C => n1609, Z => n1629);
   U1703 : OR3 port map( A => n4779, B => n4544, C => n1609, Z => n1634);
   U1707 : OR3 port map( A => n4780, B => n4543, C => n1609, Z => n1638);
   U1711 : OR3 port map( A => n4571, B => n4440, C => n1609, Z => n1642);
   U1717 : OR3 port map( A => n4387, B => n4420, C => n1609, Z => n1648);
   U1721 : OR3 port map( A => n4460, B => n4583, C => n1609, Z => n1653);
   U1725 : OR3 port map( A => n4785, B => n4415, C => n1609, Z => n1659);
   U1729 : OR3 port map( A => n4457, B => n4582, C => n1609, Z => n1663);
   U1733 : OR3 port map( A => n4788, B => n4552, C => n1609, Z => n1669);
   U1739 : OR3 port map( A => n4789, B => n4551, C => n1609, Z => n1672);
   U1747 : OR3 port map( A => n4403, B => n4570, C => n1609, Z => n1696);
   U1753 : OR3 port map( A => n4792, B => n4520, C => n1609, Z => n1699);
   U1767 : OR3 port map( A => n4388, B => n4581, C => n1609, Z => n1728);
   U1771 : OR3 port map( A => n4577, B => n4433, C => n1609, Z => n1733);
   U1775 : OR3 port map( A => n4385, B => n4580, C => n1609, Z => n1736);
   U1779 : OR3 port map( A => n4799, B => n4446, C => n1609, Z => n1740);
   U1783 : OR3 port map( A => n4576, B => n4455, C => n1609, Z => n1743);
   U1787 : OR3 port map( A => n4390, B => n4432, C => n1609, Z => n1746);
   U1791 : OR3 port map( A => n4725, B => n4445, C => n1609, Z => n1749);
   U1795 : OR3 port map( A => n4732, B => n4419, C => n1609, Z => n1752);
   U1801 : OR3 port map( A => n4575, B => n4439, C => n1609, Z => n1757);
   U1806 : OR3 port map( A => n4574, B => n4425, C => n1609, Z => n1761);
   U1811 : OR3 port map( A => n4461, B => n4618, C => n1609, Z => n1764);
   U1816 : OR3 port map( A => n4760, B => n4563, C => n1609, Z => n1768);
   U1821 : OR3 port map( A => n4761, B => n4562, C => n1609, Z => n1771);
   U1826 : OR3 port map( A => n4771, B => n4542, C => n1609, Z => n1774);
   U1831 : OR3 port map( A => n4787, B => n4617, C => n1609, Z => n1777);
   U1836 : OR3 port map( A => n4804, B => n4561, C => n1609, Z => n1781);
   U1843 : OR3 port map( A => n4459, B => n4616, C => n4352, Z => n1785);
   U1848 : OR3 port map( A => n4573, B => n4438, C => n4352, Z => n1790);
   U1853 : OR3 port map( A => n4773, B => n4510, C => n4352, Z => n1793);
   U1858 : OR3 port map( A => n4458, B => n4615, C => n4352, Z => n1796);
   U1863 : OR3 port map( A => n4572, B => n4451, C => n4352, Z => n1800);
   U1868 : OR3 port map( A => n4779, B => n4541, C => n4352, Z => n1803);
   U1873 : OR3 port map( A => n4780, B => n4560, C => n4352, Z => n1806);
   U1878 : OR3 port map( A => n4571, B => n4456, C => n4352, Z => n1809);
   U1885 : OR3 port map( A => n4387, B => n4525, C => n4352, Z => n1813);
   U1890 : OR3 port map( A => n4460, B => n4614, C => n4352, Z => n1817);
   U1895 : OR3 port map( A => n4785, B => n4524, C => n4352, Z => n1821);
   U1900 : OR3 port map( A => n4457, B => n4613, C => n4352, Z => n1824);
   U1905 : OR3 port map( A => n4788, B => n4540, C => n4352, Z => n1828);
   U1910 : OR3 port map( A => n4789, B => n4539, C => n4352, Z => n1832);
   U1915 : OR3 port map( A => n4403, B => n4568, C => n4352, Z => n1835);
   U1920 : OR3 port map( A => n4792, B => n4523, C => n4352, Z => n1839);
   U1927 : OR3 port map( A => n4388, B => n4607, C => n4352, Z => n1843);
   U1931 : OR3 port map( A => n4577, B => n4431, C => n4352, Z => n1848);
   U1935 : OR3 port map( A => n4385, B => n4606, C => n4352, Z => n1851);
   U1939 : OR3 port map( A => n4799, B => n4550, C => n4352, Z => n1855);
   U1943 : OR3 port map( A => n4576, B => n4444, C => n4352, Z => n1858);
   U1947 : OR3 port map( A => n4390, B => n4532, C => n4352, Z => n1862);
   U1957 : OR3 port map( A => n4725, B => n4605, C => n4352, Z => n1883);
   U1963 : OR3 port map( A => n4732, B => n4519, C => n4352, Z => n1887);
   U1977 : OR3 port map( A => n4459, B => n4612, C => n4706, Z => n1919);
   U1982 : OR3 port map( A => n4573, B => n4437, C => n4706, Z => n1925);
   U1987 : OR3 port map( A => n4773, B => n4611, C => n4706, Z => n1928);
   U1992 : OR3 port map( A => n4458, B => n4610, C => n4706, Z => n1932);
   U1997 : OR3 port map( A => n4572, B => n4436, C => n4706, Z => n1936);
   U2002 : OR3 port map( A => n4779, B => n4559, C => n4706, Z => n1939);
   --U2013 : AN3 port map( A => n4780, B => n4558, C => n4706, Z => n1961);--changing AN3 with OR3
   U2013 : OR3 port map( A => n4780, B => n4558, C => n4706, Z => n1961);
   --U2018 : AN3 port map( A => n4571, B => n4450, C => n4706, Z => n1964);--changing AN3 with OR3
   U2018 : OR3 port map( A => n4571, B => n4450, C => n4706, Z => n1964);
   U2028 : AN3 port map( A => v_RAM_OUT0_25_port, B => n1978, C => n4884, Z => 
                           n1974);
   U2035 : OR3 port map( A => n4387, B => n4518, C => n4706, Z => n1993);
   U2047 : OR3 port map( A => n4457, B => n4594, C => n4706, Z => n2003);
   U2051 : OR3 port map( A => n4788, B => n4531, C => n4706, Z => n2007);
   U2055 : OR3 port map( A => n4789, B => n4549, C => n4706, Z => n2010);
   U2059 : OR3 port map( A => n4403, B => n4548, C => n4706, Z => n2013);
   U2063 : OR3 port map( A => n4792, B => n4530, C => n4706, Z => n2016);
   U2070 : OR3 port map( A => n4388, B => n4418, C => n4706, Z => n2022);
   U2094 : OR3 port map( A => n4966, B => n4990, C => n4361, Z => n2077);
   U2109 : OR3 port map( A => n4577, B => n4398, C => n4706, Z => n2102);
   U2151 : OR3 port map( A => n4385, B => n4414, C => n4706, Z => n2169);
   U2186 : OR3 port map( A => n4799, B => n4566, C => n4706, Z => n2218);
   U2204 : OR3 port map( A => n4971, B => n4978, C => n4690, Z => n2237);
   U2205 : OR4 port map( A => n2241, B => n4957, C => n2243, D => n2244, Z => 
                           n2222);
   U2229 : OR3 port map( A => n4576, B => n4401, C => n4706, Z => n2267);
   U2236 : OR2 port map( A => n2032, B => n4963, Z => n2276);
   U2250 : OR2 port map( A => n2065, B => n5040, Z => n2292);
   U2271 : OR3 port map( A => n4390, B => n4430, C => n4706, Z => n2314);
   U2327 : OR3 port map( A => n4725, B => n4429, C => n4706, Z => n2351);
   U2389 : OR3 port map( A => n4732, B => n4529, C => n4706, Z => n2389);
   U2395 : OR3 port map( A => n4864, B => n2391, C => n2392, Z => n1602);
   U2526 : OR3 port map( A => n4575, B => n4435, C => n4706, Z => n2424);
   U2531 : OR3 port map( A => n4574, B => n4424, C => n4706, Z => n2428);
   U2541 : OR3 port map( A => n4760, B => n4557, C => n4706, Z => n2432);
   U2546 : OR3 port map( A => n4761, B => n4538, C => n4706, Z => n2435);
   U2553 : OR3 port map( A => n4771, B => n4537, C => n4706, Z => n2438);
   U2562 : OR3 port map( A => n4787, B => n4556, C => n4706, Z => n2461);
   U2569 : OR3 port map( A => n4804, B => n4555, C => n4706, Z => n2464);
   U2584 : OR3 port map( A => n4459, B => n4593, C => n1527, Z => n2492);
   U2596 : OR3 port map( A => n2515, B => n2516, C => n2517, Z => n2499);
   U2610 : AN3 port map( A => n2549, B => n2550, C => n5042, Z => n2548);
   U2622 : OR3 port map( A => n4573, B => n4428, C => n1527, Z => n2571);
   U2630 : AN3 port map( A => n2583, B => n2584, C => n2527, Z => n2582);
   U2656 : OR3 port map( A => n4912, B => n4901, C => n4687, Z => n2630);
   U2662 : OR3 port map( A => n4773, B => n4413, C => n1527, Z => n2637);
   U2702 : OR3 port map( A => n4458, B => n4592, C => n1527, Z => n2696);
   U2746 : OR3 port map( A => n4572, B => n4443, C => n1527, Z => n2744);
   U2793 : OR3 port map( A => n4779, B => n4528, C => n1527, Z => n2788);
   U2844 : OR3 port map( A => n4780, B => n4442, C => n1527, Z => n2825);
   U2904 : OR3 port map( A => n4571, B => n4454, C => n1527, Z => n2863);
   U2908 : OR3 port map( A => n4864, B => n2866, C => n2392, Z => n1702);
   U3037 : OR3 port map( A => n4387, B => n4522, C => n1527, Z => n2895);
   U3050 : OR3 port map( A => n2919, B => n2920, C => n2921, Z => n2901);
   U3063 : AN3 port map( A => n2953, B => n2954, C => n5037, Z => n2952);
   U3075 : OR3 port map( A => n4460, B => n4609, C => n1527, Z => n2972);
   --U3084 : OR3 port map( A => n2986, B => n2987, C => n2932, Z => n2985);--changing OR3 with AN3
   U3084 : AN3 port map( A => n2986, B => n2987, C => n2932, Z => n2985);
   U3110 : OR3 port map( A => n4935, B => n4926, C => n4682, Z => n3034);
   U3116 : OR3 port map( A => n4785, B => n4521, C => n1527, Z => n3041);
   U3157 : OR3 port map( A => n4457, B => n4608, C => n1527, Z => n3101);
   U3203 : OR3 port map( A => n4788, B => n4536, C => n1527, Z => n3148);
   U3248 : OR3 port map( A => n4789, B => n4535, C => n1527, Z => n3193);
   U3307 : OR3 port map( A => n4403, B => n4567, C => n1527, Z => n3229);
   U3368 : OR3 port map( A => n4792, B => n4534, C => n1527, Z => n3267);
   U3394 : AN3 port map( A => v_RAM_OUT0_17_port, B => n1712, C => n4938, Z => 
                           n3277);
   U3497 : OR3 port map( A => n4575, B => n4417, C => n4352, Z => n3297);
   U3509 : OR3 port map( A => n3321, B => n3322, C => n3323, Z => n3303);
   U3522 : AN3 port map( A => n3355, B => n3356, C => n5044, Z => n3354);
   U3534 : OR3 port map( A => n4574, B => n4416, C => n4352, Z => n3374);
   U3542 : AN3 port map( A => n3387, B => n3388, C => n3334, Z => n3386);
   U3568 : OR3 port map( A => n5017, B => n5008, C => n4678, Z => n3435);
   U3574 : OR3 port map( A => n4461, B => n4604, C => n4352, Z => n3442);
   U3614 : OR3 port map( A => n4760, B => n4547, C => n4352, Z => n3503);
   U3659 : OR3 port map( A => n4761, B => n4546, C => n4352, Z => n3549);
   U3703 : OR3 port map( A => n4771, B => n4517, C => n4352, Z => n3594);
   U3761 : OR3 port map( A => n4787, B => n4603, C => n4352, Z => n3630);
   U3821 : OR3 port map( A => n4804, B => n4545, C => n4352, Z => n3669);
   U3849 : AN3 port map( A => v_RAM_OUT0_1_port, B => n2476, C => n5020, Z => 
                           n3681);
   U3953 : OR3 port map( A => v_CALCULATION_CNTR_3_port, B => n4864, C => n4579
                           , Z => n3699);
   U4172 : OR2 port map( A => v_CALCULATION_CNTR_7_port, B => 
                           v_CALCULATION_CNTR_6_port, Z => n3805);
   U4178 : OR3 port map( A => v_CALCULATION_CNTR_1_port, B => n4864, C => n4384
                           , Z => n3800);
   U4199 : OR3 port map( A => v_CALCULATION_CNTR_5_port, B => 
                           v_CALCULATION_CNTR_7_port, C => 
                           v_CALCULATION_CNTR_6_port, Z => n3809);
   U104 : EOI port map( A => n116, B => n117, Z => n115);
   U105 : EOI port map( A => n118, B => n119, Z => n117);
   U106 : EOI port map( A => n120, B => n121, Z => n116);
   U107 : EOI port map( A => n122, B => n123, Z => n113);
   U108 : EOI port map( A => n124, B => n125, Z => n123);
   U109 : EOI port map( A => n126, B => n127, Z => n122);
   U110 : EOI port map( A => n128, B => n129, Z => n109);
   U111 : EOI port map( A => n130, B => n131, Z => n129);
   --U112 : EOI port map( A => n132, B => n133, Z => n128);--changing EOI with ENI
   U112 : ENI port map( A => n132, B => n133, Z => n128);
   U114 : EOI port map( A => n138, B => n139, Z => n136);
   U115 : EOI port map( A => n140, B => n141, Z => n139);
   U116 : ENI port map( A => n142, B => n143, Z => n138);
   U117 : EOI port map( A => v_KEY_COLUMN_9_port, B => v_DATA_COLUMN_9_port, Z 
                           => n135);
   U119 : AO1P port map( A => n147, B => n4386, C => n149, D => n150, Z => n146
                           );
   U120 : NR2I port map( A => n4383, B => n151, Z => n150);
   -- U121 : NR2I port map( A => n152, B => n153, Z => n151);--changing NR2I with EOI
   U121 : EOI port map( A => n152, B => n153, Z => n151);
   U122 : EOI port map( A => n154, B => n155, Z => n153);
   U123 : EOI port map( A => n156, B => n157, Z => n155);
   U124 : EOI port map( A => n158, B => n159, Z => n152);
   U125 : EOI port map( A => n160, B => n161, Z => n159);
   U127 : EOI port map( A => n166, B => n167, Z => n165);
   U128 : EOI port map( A => n168, B => n169, Z => n167);
   U129 : EOI port map( A => n170, B => n171, Z => n169);
   U130 : EOI port map( A => n172, B => n173, Z => n166);
   U131 : EOI port map( A => n174, B => n175, Z => n173);
   U132 : EOI port map( A => v_DATA_COLUMN_8_port, B => n4732, Z => n162);
   U133 : EOI port map( A => n177, B => n178, Z => n147);
   U134 : EOI port map( A => n179, B => n180, Z => n178);
   U135 : EOI port map( A => n181, B => n182, Z => n180);
   U136 : EOI port map( A => n183, B => n184, Z => n177);
   U137 : ENI port map( A => n185, B => n186, Z => n183);
   U144 : EOI port map( A => n4807, B => n201_port, Z => n192_port);
   U148 : ENI port map( A => n203_port, B => n204, Z => n196);
   --U152 : ENI port map( A => n212, B => n213, Z => n211);--changing ENI with EOI
   U152 : EOI port map( A => n212, B => n213, Z => n211);
   U153 : ENI port map( A => n214, B => n215, Z => n213);
   U154 : EOI port map( A => n160, B => n216, Z => n212);
   U155 : EOI port map( A => n217, B => n218, Z => n210);
   U156 : ENI port map( A => n219, B => n220, Z => n218);
   U157 : EOI port map( A => n181, B => n221, Z => n217);
   U158 : EOI port map( A => n222, B => n223, Z => n208);
   U159 : EOI port map( A => n174, B => n224, Z => n223);
   U160 : EOI port map( A => n225, B => n226, Z => n222);
   U162 : EOI port map( A => n229, B => n230, Z => n228);
   U163 : EOI port map( A => n204, B => n231, Z => n230);
   U164 : ENI port map( A => n232, B => n233, Z => n229);
   U165 : EOI port map( A => n4657, B => v_DATA_COLUMN_7_port, Z => n227);
   U169 : EOI port map( A => n241, B => n242, Z => n240);
   U170 : EOI port map( A => n243, B => n244, Z => n241);
   U171 : EOI port map( A => n245, B => n246, Z => n239);
   U172 : EOI port map( A => n247, B => n248, Z => n245);
   U173 : EOI port map( A => n249, B => n250, Z => n237);
   U174 : EOI port map( A => n251, B => n252, Z => n250);
   U176 : EOI port map( A => n255, B => n256, Z => n254);
   U177 : EOI port map( A => n257, B => n258, Z => n255);
   U178 : EOI port map( A => n4656, B => v_DATA_COLUMN_6_port, Z => n253);
   U182 : EOI port map( A => n266, B => n267, Z => n265);
   U183 : EOI port map( A => n268, B => n269, Z => n267);
   U184 : EOI port map( A => n270, B => n271, Z => n266);
   U185 : EOI port map( A => n272, B => n273, Z => n264);
   U186 : EOI port map( A => n274, B => n275, Z => n273);
   U187 : EOI port map( A => n276, B => n277, Z => n272);
   U188 : EOI port map( A => n278, B => n279, Z => n262);
   U189 : EOI port map( A => n280, B => n281, Z => n279);
   U190 : ENI port map( A => n282, B => n283, Z => n278);
   U192 : EOI port map( A => n286, B => n287, Z => n285);
   U193 : EOI port map( A => n288, B => n289, Z => n287);
   U194 : ENI port map( A => n290, B => n291, Z => n286);
   U195 : EOI port map( A => n4655, B => v_DATA_COLUMN_5_port, Z => n284);
   U199 : EOI port map( A => n299, B => n300, Z => n298);
   U200 : EOI port map( A => n301, B => n302, Z => n300);
   U201 : EOI port map( A => n303, B => n304, Z => n299);
   U202 : EOI port map( A => n305, B => n306, Z => n297);
   U203 : EOI port map( A => n307, B => n308, Z => n306);
   U204 : EOI port map( A => n309, B => n310, Z => n305);
   U205 : EOI port map( A => n311, B => n312, Z => n295);
   U206 : EOI port map( A => n313, B => n314, Z => n312);
   U207 : EOI port map( A => n315, B => n316, Z => n311);
   U209 : EOI port map( A => n319, B => n320, Z => n318);
   U210 : EOI port map( A => n321, B => n322, Z => n320);
   U211 : EOI port map( A => n323, B => n324, Z => n319);
   U212 : EOI port map( A => v_KEY_COLUMN_4_port, B => v_DATA_COLUMN_4_port, Z 
                           => n317);
   U216 : EOI port map( A => n332, B => n333, Z => n331);
   U217 : EOI port map( A => n334, B => n335, Z => n333);
   U218 : EOI port map( A => n336, B => n337, Z => n332);
   U219 : EOI port map( A => n338, B => n339, Z => n337);
   U220 : EOI port map( A => n340, B => n341, Z => n330);
   U221 : EOI port map( A => n342, B => n343, Z => n341);
   U222 : EOI port map( A => n344, B => n345, Z => n340);
   U223 : EOI port map( A => n346, B => n347, Z => n345);
   U224 : EOI port map( A => n348, B => n349, Z => n328);
   U225 : EOI port map( A => n350, B => n351, Z => n349);
   U226 : EOI port map( A => n352, B => n353, Z => n351);
   U227 : ENI port map( A => n354, B => n355, Z => n348);
   U229 : EOI port map( A => n358, B => n359, Z => n357);
   U230 : EOI port map( A => n360, B => n361, Z => n359);
   U231 : EOI port map( A => n362, B => n363, Z => n361);
   U232 : ENI port map( A => n364, B => n365, Z => n358);
   U233 : EOI port map( A => v_KEY_COLUMN_3_port, B => v_DATA_COLUMN_3_port, Z 
                           => n356);
   U237 : EOI port map( A => n373, B => n374, Z => n372);
   U238 : EOI port map( A => n161, B => n375, Z => n373);
   U239 : EOI port map( A => n376, B => n216, Z => n375);
   U240 : EOI port map( A => n377, B => n378, Z => n371);
   U241 : EOI port map( A => n182, B => n379, Z => n377);
   U242 : EOI port map( A => n380, B => n221, Z => n379);
   U243 : EOI port map( A => n381, B => n382, Z => n369);
   U244 : EOI port map( A => n175, B => n383, Z => n382);
   U245 : EOI port map( A => n384, B => n224, Z => n383);
   U247 : EOI port map( A => n387, B => n388, Z => n386);
   U248 : EOI port map( A => n231, B => n389, Z => n388);
   U249 : EOI port map( A => n203_port, B => n390, Z => n389);
   U250 : EOI port map( A => n4671, B => v_DATA_COLUMN_31_port, Z => n385);
   U254 : EOI port map( A => n398, B => n399, Z => n397);
   U255 : EOI port map( A => n400, B => n401, Z => n398);
   U256 : EOI port map( A => n402, B => n403, Z => n401);
   U257 : EOI port map( A => n404, B => n405, Z => n396);
   U258 : EOI port map( A => n406, B => n407, Z => n404);
   U259 : EOI port map( A => n408, B => n409, Z => n407);
   U260 : EOI port map( A => n410, B => n411, Z => n394);
   U261 : EOI port map( A => n412, B => n413, Z => n411);
   U262 : EOI port map( A => n414, B => n415, Z => n413);
   U264 : EOI port map( A => n418, B => n419, Z => n417);
   U265 : EOI port map( A => n420, B => n421, Z => n419);
   U266 : EOI port map( A => n422, B => n423, Z => n421);
   U267 : EOI port map( A => n4670, B => v_DATA_COLUMN_30_port, Z => n416);
   U271 : EOI port map( A => n431, B => n432, Z => n430);
   U272 : EOI port map( A => n433, B => n434, Z => n432);
   U273 : ENI port map( A => n435, B => n436, Z => n431);
   U274 : ENI port map( A => n437, B => n438, Z => n436);
   U275 : EOI port map( A => n439, B => n440, Z => n429);
   U276 : EOI port map( A => n441, B => n442, Z => n440);
   U277 : ENI port map( A => n443, B => n444, Z => n439);
   U278 : ENI port map( A => n445, B => n446, Z => n444);
   U279 : EOI port map( A => n447, B => n448, Z => n427);
   U280 : EOI port map( A => n449, B => n450, Z => n448);
   U281 : ENI port map( A => n451, B => n452, Z => n450);
   U282 : ENI port map( A => n453, B => n454, Z => n447);
   U284 : EOI port map( A => n457, B => n458, Z => n456);
   U285 : EOI port map( A => n459, B => n460, Z => n458);
   U286 : EOI port map( A => n461, B => n462, Z => n460);
   U287 : ENI port map( A => n463, B => n464, Z => n457);
   U288 : EOI port map( A => v_KEY_COLUMN_2_port, B => v_DATA_COLUMN_2_port, Z 
                           => n455);
   U292 : EOI port map( A => n472, B => n473, Z => n471);
   U293 : EOI port map( A => n269, B => n474, Z => n473);
   U294 : EOI port map( A => n475, B => n476, Z => n269);
   U295 : EOI port map( A => n243, B => n477, Z => n472);
   U296 : EOI port map( A => n478, B => n479, Z => n470);
   U297 : EOI port map( A => n275, B => n480, Z => n479);
   U298 : EOI port map( A => n481, B => n482, Z => n275);
   U299 : EOI port map( A => n247, B => n483, Z => n478);
   U300 : EOI port map( A => n484, B => n485, Z => n468);
   U301 : EOI port map( A => n251, B => n486, Z => n485);
   U302 : EOI port map( A => n487, B => n282, Z => n484);
   U303 : EOI port map( A => n488, B => n489, Z => n282);
   U305 : EOI port map( A => n492, B => n493, Z => n491);
   U306 : EOI port map( A => n258, B => n494, Z => n493);
   U307 : EOI port map( A => n495, B => n290, Z => n492);
   U308 : EOI port map( A => n496, B => n497, Z => n290);
   U309 : EOI port map( A => v_KEY_COLUMN_29_port, B => v_DATA_COLUMN_29_port, 
                           Z => n490);
   U313 : EOI port map( A => n505, B => n506, Z => n504);
   U314 : EOI port map( A => n507, B => n508, Z => n506);
   U315 : EOI port map( A => n271, B => n304, Z => n505);
   U316 : EOI port map( A => n509, B => n510, Z => n503);
   U317 : EOI port map( A => n511, B => n512, Z => n510);
   U318 : EOI port map( A => n277, B => n310, Z => n509);
   U319 : EOI port map( A => n513, B => n514, Z => n501);
   U320 : EOI port map( A => n281, B => n314, Z => n514);
   U321 : EOI port map( A => n515, B => n516, Z => n513);
   U323 : EOI port map( A => n519, B => n520, Z => n518);
   U324 : EOI port map( A => n289, B => n322, Z => n520);
   U325 : EOI port map( A => n521, B => n522, Z => n519);
   U326 : EOI port map( A => n4669, B => v_DATA_COLUMN_28_port, Z => n517);
   U330 : EOI port map( A => n530, B => n531, Z => n529);
   U331 : EOI port map( A => n532, B => n533, Z => n531);
   U332 : EOI port map( A => n534, B => n535, Z => n530);
   U333 : EOI port map( A => n536, B => n339, Z => n535);
   U334 : EOI port map( A => n537, B => n538, Z => n528);
   U335 : EOI port map( A => n539, B => n540, Z => n538);
   U336 : EOI port map( A => n541, B => n542, Z => n537);
   U337 : EOI port map( A => n543, B => n347, Z => n542);
   U338 : EOI port map( A => n544, B => n545, Z => n526);
   U339 : EOI port map( A => n546, B => n547, Z => n545);
   U340 : EOI port map( A => n548, B => n353, Z => n547);
   U341 : EOI port map( A => n549, B => n4730, Z => n544);
   U344 : EOI port map( A => n554, B => n555, Z => n553);
   U345 : EOI port map( A => n360, B => n556, Z => n555);
   U346 : EOI port map( A => n557, B => n558, Z => n556);
   U347 : EOI port map( A => n559, B => n4729, Z => n554);
   U349 : EOI port map( A => n4668, B => v_DATA_COLUMN_27_port, Z => n552);
   U353 : EOI port map( A => n569, B => n570, Z => n568);
   U354 : EOI port map( A => n571, B => n572, Z => n570);
   U355 : EOI port map( A => n573, B => n574, Z => n569);
   U356 : EOI port map( A => n575, B => n576, Z => n567);
   U357 : EOI port map( A => n577, B => n578, Z => n576);
   U358 : EOI port map( A => n579, B => n580, Z => n575);
   U359 : EOI port map( A => n581, B => n582, Z => n565);
   U360 : EOI port map( A => n583, B => n584, Z => n582);
   U361 : EOI port map( A => n585, B => n586, Z => n581);
   U363 : EOI port map( A => n589, B => n590, Z => n588);
   U364 : EOI port map( A => n591, B => n592, Z => n590);
   U365 : EOI port map( A => n593, B => n594, Z => n589);
   U366 : EOI port map( A => v_KEY_COLUMN_26_port, B => v_DATA_COLUMN_26_port, 
                           Z => n587);
   U370 : EOI port map( A => n602, B => n603, Z => n601);
   U371 : EOI port map( A => n604, B => n605, Z => n603);
   U372 : ENI port map( A => n118, B => n437, Z => n602);
   U373 : EOI port map( A => n606, B => n607, Z => n600);
   U374 : EOI port map( A => n608, B => n609, Z => n607);
   U375 : ENI port map( A => n124, B => n445, Z => n606);
   U376 : EOI port map( A => n610, B => n611, Z => n598);
   U377 : ENI port map( A => n133, B => n451, Z => n611);
   U378 : EOI port map( A => n612, B => n4762, Z => n610);
   U380 : EOI port map( A => n616, B => n617, Z => n615);
   U381 : EOI port map( A => n140, B => n461, Z => n617);
   U382 : EOI port map( A => n618, B => n4763, Z => n616);
   U383 : EOI port map( A => v_KEY_COLUMN_25_port, B => v_DATA_COLUMN_25_port, 
                           Z => n614);
   U387 : EOI port map( A => n627, B => n628, Z => n626);
   U388 : EOI port map( A => n629, B => n630, Z => n628);
   U389 : EOI port map( A => n154, B => n631, Z => n630);
   U390 : EOI port map( A => n157, B => n632, Z => n627);
   U391 : EOI port map( A => n633, B => n634, Z => n632);
   U392 : EOI port map( A => n635, B => n636, Z => n625);
   U393 : EOI port map( A => n4731, B => n638, Z => n636);
   U394 : EOI port map( A => n184, B => n639, Z => n638);
   U396 : EOI port map( A => n185, B => n641, Z => n635);
   U397 : EOI port map( A => n642, B => n643, Z => n641);
   U398 : EOI port map( A => n644, B => n645, Z => n623);
   U399 : EOI port map( A => n171, B => n646, Z => n645);
   U400 : EOI port map( A => n647, B => n648, Z => n646);
   U401 : EOI port map( A => n649, B => n650, Z => n644);
   U402 : EOI port map( A => n4738, B => n168, Z => n649);
   U404 : EOI port map( A => n654, B => n655, Z => n653);
   U405 : EOI port map( A => n656, B => n657, Z => n655);
   U406 : EOI port map( A => n658, B => n659, Z => n657);
   U407 : EOI port map( A => n660, B => n661, Z => n654);
   U408 : EOI port map( A => n4742, B => n201_port, Z => n660);
   U409 : EOI port map( A => n4667, B => v_DATA_COLUMN_24_port, Z => n652);
   U413 : EOI port map( A => n670, B => n374, Z => n669);
   U414 : EOI port map( A => n671, B => n672, Z => n374);
   U415 : EOI port map( A => n673, B => n674, Z => n672);
   U416 : ENI port map( A => n214, B => n675, Z => n670);
   U417 : EOI port map( A => n633, B => n676, Z => n675);
   U418 : EOI port map( A => n677, B => n378, Z => n668);
   U419 : EOI port map( A => n678, B => n679, Z => n378);
   U420 : EOI port map( A => n680, B => n681, Z => n679);
   U421 : ENI port map( A => n219, B => n682, Z => n677);
   U422 : EOI port map( A => n642, B => n683, Z => n682);
   U423 : EOI port map( A => n381, B => n684, Z => n666);
   U424 : EOI port map( A => n4753, B => n686, Z => n684);
   U425 : EOI port map( A => n647, B => n687, Z => n686);
   U426 : EOI port map( A => n688, B => n689, Z => n381);
   U427 : EOI port map( A => n4768, B => n691, Z => n688);
   U429 : EOI port map( A => n387, B => n694, Z => n693);
   U430 : EOI port map( A => n233, B => n695, Z => n694);
   U431 : EOI port map( A => n658, B => n696, Z => n695);
   U432 : EOI port map( A => n697, B => n4741, Z => n387);
   U433 : EOI port map( A => n4769, B => n700, Z => n697);
   U434 : EOI port map( A => n4666, B => v_DATA_COLUMN_23_port, Z => n692);
   U438 : EOI port map( A => n708, B => n242, Z => n707);
   U439 : EOI port map( A => n709, B => n710, Z => n242);
   U440 : ENI port map( A => n711, B => n154, Z => n709);
   U441 : EOI port map( A => n216, B => n712, Z => n708);
   U442 : EOI port map( A => n400, B => n270, Z => n712);
   U443 : EOI port map( A => n713, B => n246, Z => n706);
   U444 : EOI port map( A => n714, B => n715, Z => n246);
   U445 : ENI port map( A => n716, B => n184, Z => n714);
   U446 : EOI port map( A => n221, B => n717, Z => n713);
   U447 : EOI port map( A => n406, B => n276, Z => n717);
   U448 : EOI port map( A => n249, B => n718, Z => n704);
   U449 : EOI port map( A => n224, B => n719, Z => n718);
   U450 : EOI port map( A => n412, B => n280, Z => n719);
   U451 : EOI port map( A => n720, B => n721, Z => n249);
   U452 : EOI port map( A => n722, B => n168, Z => n720);
   U454 : EOI port map( A => n725, B => n726, Z => n724);
   U455 : EOI port map( A => n420, B => n288, Z => n726);
   U456 : EOI port map( A => n257, B => n231, Z => n725);
   U457 : EOI port map( A => n727, B => n728, Z => n257);
   U458 : EOI port map( A => n729, B => n201_port, Z => n727);
   U459 : EOI port map( A => n4665, B => v_DATA_COLUMN_22_port, Z => n723);
   U463 : EOI port map( A => n737, B => n738, Z => n736);
   U464 : EOI port map( A => n268, B => n475, Z => n738);
   U465 : EOI port map( A => n376, B => n739, Z => n268);
   U466 : EOI port map( A => n303, B => n740, Z => n737);
   U467 : EOI port map( A => n403, B => n477, Z => n740);
   U468 : EOI port map( A => n741, B => n742, Z => n735);
   U469 : EOI port map( A => n274, B => n481, Z => n742);
   U470 : EOI port map( A => n380, B => n743, Z => n274);
   U471 : EOI port map( A => n309, B => n744, Z => n741);
   U472 : EOI port map( A => n409, B => n483, Z => n744);
   U473 : EOI port map( A => n745, B => n746, Z => n733);
   U474 : EOI port map( A => n313, B => n747, Z => n746);
   U475 : EOI port map( A => n415, B => n486, Z => n747);
   U476 : ENI port map( A => n488, B => n283, Z => n745);
   U477 : EOI port map( A => n384, B => n748, Z => n283);
   U479 : EOI port map( A => n751, B => n752, Z => n750);
   U480 : EOI port map( A => n494, B => n753, Z => n752);
   U481 : EOI port map( A => n423, B => n321, Z => n753);
   U482 : ENI port map( A => n496, B => n291, Z => n751);
   U483 : EOI port map( A => n390, B => n754, Z => n291);
   U484 : EOI port map( A => v_KEY_COLUMN_21_port, B => v_DATA_COLUMN_21_port, 
                           Z => n749);
   U488 : EOI port map( A => n762, B => n763, Z => n761);
   U489 : EOI port map( A => n507, B => n302, Z => n763);
   U490 : ENI port map( A => n764, B => n765, Z => n302);
   U491 : EOI port map( A => n766, B => n767, Z => n764);
   U492 : EOI port map( A => n476, B => n768, Z => n762);
   U493 : EOI port map( A => n769, B => n770, Z => n760);
   U494 : EOI port map( A => n511, B => n308, Z => n770);
   U495 : ENI port map( A => n771, B => n772, Z => n308);
   U496 : EOI port map( A => n773, B => n774, Z => n771);
   U497 : EOI port map( A => n482, B => n775, Z => n769);
   U498 : EOI port map( A => n776, B => n777, Z => n758);
   U499 : EOI port map( A => n489, B => n778, Z => n777);
   U500 : EOI port map( A => n315, B => n516, Z => n776);
   U501 : EOI port map( A => n779, B => n780, Z => n315);
   U502 : EOI port map( A => n781, B => n782, Z => n779);
   U504 : EOI port map( A => n785, B => n786, Z => n784);
   U505 : EOI port map( A => n497, B => n787, Z => n786);
   U506 : EOI port map( A => n323, B => n522, Z => n785);
   U507 : EOI port map( A => n788, B => n789, Z => n323);
   U508 : EOI port map( A => n790, B => n4774, Z => n788);
   U509 : EOI port map( A => n4664, B => v_DATA_COLUMN_20_port, Z => n783);
   U513 : EOI port map( A => n799, B => n800, Z => n798);
   U514 : EOI port map( A => n801, B => n605, Z => n800);
   U515 : ENI port map( A => n802, B => n803, Z => n605);
   U516 : ENI port map( A => n804, B => n805, Z => n802);
   U517 : EOI port map( A => n120, B => n806, Z => n799);
   U518 : EOI port map( A => n807, B => n808, Z => n797);
   U519 : EOI port map( A => n809, B => n609, Z => n808);
   U520 : ENI port map( A => n810, B => n811, Z => n609);
   U521 : ENI port map( A => n812, B => n813, Z => n810);
   U522 : EOI port map( A => n126, B => n814, Z => n807);
   U523 : EOI port map( A => n815, B => n816, Z => n795);
   U524 : EOI port map( A => n130, B => n817, Z => n816);
   U525 : EOI port map( A => n612, B => n818, Z => n815);
   U526 : EOI port map( A => n819, B => n820, Z => n612);
   U527 : ENI port map( A => n821, B => n822, Z => n819);
   U529 : EOI port map( A => n825, B => n826, Z => n824);
   U530 : EOI port map( A => n141, B => n827, Z => n826);
   U531 : EOI port map( A => n618, B => n828, Z => n825);
   U532 : EOI port map( A => n829, B => n4727, Z => n618);
   U534 : ENI port map( A => n832, B => n833, Z => n829);
   U535 : EOI port map( A => v_KEY_COLUMN_1_port, B => v_DATA_COLUMN_1_port, Z 
                           => n823);
   U539 : EOI port map( A => n841, B => n842, Z => n840);
   U540 : EOI port map( A => n334, B => n532, Z => n842);
   U541 : ENI port map( A => n843, B => n844, Z => n532);
   U542 : EOI port map( A => n4800, B => n846, Z => n843);
   U543 : ENI port map( A => n847, B => n848, Z => n334);
   U544 : EOI port map( A => n534, B => n849, Z => n841);
   U545 : EOI port map( A => n850, B => n851, Z => n849);
   U546 : EOI port map( A => n852, B => n853, Z => n839);
   U547 : EOI port map( A => n342, B => n539, Z => n853);
   U548 : ENI port map( A => n854, B => n855, Z => n539);
   U549 : EOI port map( A => n4801, B => n857, Z => n854);
   U550 : ENI port map( A => n858, B => n859, Z => n342);
   U551 : EOI port map( A => n541, B => n860, Z => n852);
   U552 : EOI port map( A => n861, B => n862, Z => n860);
   U553 : EOI port map( A => n863, B => n864, Z => n837);
   U554 : EOI port map( A => n546, B => n865, Z => n864);
   U555 : EOI port map( A => n866, B => n867, Z => n865);
   U556 : EOI port map( A => n551, B => n355, Z => n863);
   U557 : ENI port map( A => n868, B => n869, Z => n355);
   U558 : EOI port map( A => n870, B => n871, Z => n551);
   U559 : EOI port map( A => n4802, B => n873, Z => n870);
   U561 : EOI port map( A => n876, B => n877, Z => n875);
   U562 : EOI port map( A => n878, B => n879, Z => n877);
   U563 : EOI port map( A => n880, B => n558, Z => n879);
   U564 : EOI port map( A => n559, B => n364, Z => n876);
   U565 : EOI port map( A => n881, B => n882, Z => n364);
   U566 : EOI port map( A => n883, B => n884, Z => n559);
   U567 : EOI port map( A => n4803, B => n886, Z => n883);
   U568 : EOI port map( A => v_KEY_COLUMN_19_port, B => v_DATA_COLUMN_19_port, 
                           Z => n874);
   U572 : EOI port map( A => n894, B => n895, Z => n893);
   U573 : EOI port map( A => n433, B => n572, Z => n895);
   U574 : ENI port map( A => n896, B => n897, Z => n572);
   U575 : ENI port map( A => n438, B => n898, Z => n896);
   U576 : EOI port map( A => n899, B => n804, Z => n433);
   U577 : EOI port map( A => n900, B => n901, Z => n894);
   U578 : EOI port map( A => n121, B => n806, Z => n901);
   U579 : EOI port map( A => n902, B => n903, Z => n892);
   U580 : EOI port map( A => n441, B => n578, Z => n903);
   U581 : ENI port map( A => n904, B => n905, Z => n578);
   U582 : ENI port map( A => n446, B => n906, Z => n904);
   U583 : EOI port map( A => n907, B => n812, Z => n441);
   U584 : EOI port map( A => n908, B => n909, Z => n902);
   U585 : EOI port map( A => n127, B => n814, Z => n909);
   U586 : EOI port map( A => n910, B => n911, Z => n890);
   U587 : EOI port map( A => n912, B => n913, Z => n911);
   U588 : EOI port map( A => n131, B => n817, Z => n913);
   U589 : EOI port map( A => n585, B => n454, Z => n910);
   U590 : EOI port map( A => n914, B => n821, Z => n454);
   U591 : EOI port map( A => n915, B => n916, Z => n585);
   U592 : ENI port map( A => n452, B => n917, Z => n915);
   U594 : EOI port map( A => n920, B => n921, Z => n919);
   U595 : EOI port map( A => n922, B => n923, Z => n921);
   U596 : EOI port map( A => n143, B => n827, Z => n923);
   U597 : EOI port map( A => n593, B => n463, Z => n920);
   U598 : EOI port map( A => n832, B => n924, Z => n463);
   U599 : EOI port map( A => n925, B => n926, Z => n593);
   U600 : EOI port map( A => n4772, B => n462, Z => n925);
   U602 : EOI port map( A => v_KEY_COLUMN_18_port, B => v_DATA_COLUMN_18_port, 
                           Z => n918);
   U606 : EOI port map( A => n936, B => n937, Z => n935);
   U607 : EOI port map( A => n604, B => n801, Z => n937);
   U608 : ENI port map( A => n119, B => n435, Z => n936);
   U609 : ENI port map( A => n938, B => n573, Z => n119);
   U610 : ENI port map( A => n437, B => n806, Z => n573);
   U611 : ENI port map( A => n899, B => n805, Z => n938);
   U612 : ENI port map( A => n939, B => n940, Z => n805);
   U613 : EOI port map( A => n154, B => n244, Z => n940);
   U614 : EOI port map( A => n676, B => n403, Z => n244);
   U615 : EOI port map( A => n941, B => n216, Z => n939);
   U616 : ENI port map( A => n270, B => n376, Z => n941);
   U617 : EOI port map( A => n942, B => n943, Z => n934);
   U618 : EOI port map( A => n608, B => n809, Z => n943);
   U619 : ENI port map( A => n125, B => n443, Z => n942);
   U620 : ENI port map( A => n944, B => n579, Z => n125);
   U621 : ENI port map( A => n445, B => n814, Z => n579);
   U622 : ENI port map( A => n907, B => n813, Z => n944);
   U623 : ENI port map( A => n945, B => n946, Z => n813);
   U624 : EOI port map( A => n184, B => n248, Z => n946);
   U625 : EOI port map( A => n683, B => n409, Z => n248);
   U626 : EOI port map( A => n947, B => n221, Z => n945);
   U627 : ENI port map( A => n276, B => n380, Z => n947);
   U628 : EOI port map( A => n948, B => n949, Z => n932);
   U629 : EOI port map( A => n132, B => n449, Z => n949);
   U630 : ENI port map( A => n950, B => n583, Z => n132);
   U631 : ENI port map( A => n451, B => n817, Z => n583);
   U632 : ENI port map( A => n914, B => n822, Z => n950);
   U633 : ENI port map( A => n951, B => n952, Z => n822);
   U634 : EOI port map( A => n168, B => n252, Z => n952);
   U635 : EOI port map( A => n687, B => n415, Z => n252);
   U636 : EOI port map( A => n953, B => n224, Z => n951);
   U637 : ENI port map( A => n280, B => n384, Z => n953);
   U638 : EOI port map( A => n954, B => n818, Z => n948);
   U640 : EOI port map( A => n957, B => n958, Z => n956);
   U641 : EOI port map( A => n142, B => n459, Z => n958);
   U642 : ENI port map( A => n959, B => n591, Z => n142);
   U643 : EOI port map( A => n827, B => n461, Z => n591);
   U644 : ENI port map( A => n833, B => n924, Z => n959);
   U645 : ENI port map( A => n960, B => n961, Z => n833);
   U646 : EOI port map( A => n201_port, B => n256, Z => n961);
   U647 : EOI port map( A => n696, B => n423, Z => n256);
   U648 : EOI port map( A => n962, B => n231, Z => n960);
   U649 : EOI port map( A => n4786, B => n390, Z => n962);
   U650 : EOI port map( A => n964, B => n828, Z => n957);
   U651 : EOI port map( A => n4663, B => v_DATA_COLUMN_17_port, Z => n955);
   U653 : AO1P port map( A => n968, B => n4386, C => n969, D => n970, Z => n967
                           );
   U654 : NR2I port map( A => n4383, B => n971, Z => n970);
   U655 : EOI port map( A => n972, B => n973, Z => n971);
   U656 : EOI port map( A => n974, B => n975, Z => n973);
   U657 : EOI port map( A => n157, B => n976, Z => n972);
   U658 : EOI port map( A => n977, B => n156, Z => n976);
   U660 : EOI port map( A => n980, B => n981, Z => n979);
   U661 : EOI port map( A => n982, B => n983, Z => n981);
   U662 : EOI port map( A => n171, B => n984, Z => n980);
   U663 : EOI port map( A => n985, B => n170, Z => n984);
   U664 : EOI port map( A => v_DATA_COLUMN_16_port, B => n4792, Z => n978);
   U665 : EOI port map( A => n987, B => n988, Z => n968);
   U666 : EOI port map( A => n185, B => n989, Z => n988);
   U667 : EOI port map( A => n990, B => n186, Z => n989);
   U668 : ENI port map( A => n991, B => n992, Z => n987);
   U677 : ENI port map( A => n4807, B => n4751, Z => n1003);
   U682 : EOI port map( A => n1013, B => n1014, Z => n1012);
   U683 : EOI port map( A => n215, B => n631, Z => n1014);
   U684 : ENI port map( A => n1015, B => n674, Z => n215);
   U685 : ENI port map( A => n711, B => n767, Z => n674);
   U686 : EOI port map( A => n4795, B => n974, Z => n1015);
   U687 : EOI port map( A => n161, B => n633, Z => n974);
   U688 : EOI port map( A => n676, B => n376, Z => n1013);
   U689 : EOI port map( A => n1017, B => n1018, Z => n1011);
   U690 : EOI port map( A => n220, B => n639, Z => n1018);
   U691 : ENI port map( A => n1019, B => n681, Z => n220);
   U692 : ENI port map( A => n716, B => n774, Z => n681);
   U693 : EOI port map( A => n4796, B => n991, Z => n1019);
   U694 : ENI port map( A => n4783, B => n642, Z => n991);
   U695 : EOI port map( A => n683, B => n380, Z => n1017);
   U696 : EOI port map( A => n1022, B => n1023, Z => n1009);
   U697 : EOI port map( A => n687, B => n384, Z => n1023);
   U698 : EOI port map( A => n4738, B => n225, Z => n1022);
   U699 : ENI port map( A => n1024, B => n691, Z => n225);
   U700 : EOI port map( A => n4758, B => n782, Z => n691);
   U701 : EOI port map( A => n4797, B => n982, Z => n1024);
   U702 : EOI port map( A => n175, B => n647, Z => n982);
   U705 : EOI port map( A => n1029, B => n1030, Z => n1028);
   U706 : EOI port map( A => n696, B => n390, Z => n1030);
   U707 : EOI port map( A => n4742, B => n232, Z => n1029);
   U708 : ENI port map( A => n1031, B => n700, Z => n232);
   U709 : EOI port map( A => n4759, B => n4774, Z => n700);
   U711 : EOI port map( A => n4798, B => n4765, Z => n1031);
   U713 : ENI port map( A => n203_port, B => n658, Z => n998);
   U715 : EOI port map( A => n4662, B => v_DATA_COLUMN_15_port, Z => n1027);
   U719 : EOI port map( A => n1042, B => n399, Z => n1041);
   U720 : EOI port map( A => n710, B => n1043, Z => n399);
   U721 : EOI port map( A => n767, B => n975, Z => n1043);
   U722 : EOI port map( A => n271, B => n477, Z => n767);
   U723 : EOI port map( A => n1044, B => n739, Z => n710);
   U724 : EOI port map( A => n768, B => n304, Z => n739);
   U725 : ENI port map( A => n846, B => n4736, Z => n304);
   U726 : EOI port map( A => n270, B => n1046, Z => n1042);
   U727 : EOI port map( A => n673, B => n243, Z => n1046);
   U728 : EOI port map( A => n1047, B => n405, Z => n1040);
   U729 : EOI port map( A => n715, B => n1048, Z => n405);
   U730 : EOI port map( A => n774, B => n992, Z => n1048);
   U731 : EOI port map( A => n277, B => n483, Z => n774);
   U732 : EOI port map( A => n1049, B => n743, Z => n715);
   U733 : EOI port map( A => n775, B => n310, Z => n743);
   U734 : ENI port map( A => n857, B => n4740, Z => n310);
   U735 : EOI port map( A => n276, B => n1051, Z => n1047);
   U736 : EOI port map( A => n680, B => n247, Z => n1051);
   U737 : EOI port map( A => n410, B => n1052, Z => n1038);
   U738 : EOI port map( A => n280, B => n1053, Z => n1052);
   U739 : EOI port map( A => n1054, B => n251, Z => n1053);
   U740 : EOI port map( A => n1055, B => n721, Z => n410);
   U741 : EOI port map( A => n1056, B => n748, Z => n721);
   U742 : EOI port map( A => n778, B => n314, Z => n748);
   U743 : ENI port map( A => n873, B => n4738, Z => n314);
   U744 : ENI port map( A => n782, B => n983, Z => n1055);
   U745 : EOI port map( A => n281, B => n486, Z => n782);
   U747 : EOI port map( A => n418, B => n1059, Z => n1058);
   U748 : EOI port map( A => n288, B => n1060, Z => n1059);
   U749 : EOI port map( A => n1061, B => n258, Z => n1060);
   U750 : EOI port map( A => n1062, B => n728, Z => n418);
   U751 : EOI port map( A => n1063, B => n754, Z => n728);
   U752 : EOI port map( A => n787, B => n322, Z => n754);
   U753 : ENI port map( A => n886, B => n4742, Z => n322);
   U754 : EOI port map( A => n1033, B => n4751, Z => n1062);
   U755 : ENI port map( A => n289, B => n494, Z => n1033);
   U756 : EOI port map( A => n4661, B => v_DATA_COLUMN_14_port, Z => n1057);
   U760 : EOI port map( A => n1071, B => n1072, Z => n1070);
   U761 : EOI port map( A => n475, B => n474, Z => n1072);
   U762 : ENI port map( A => n214, B => n1044, Z => n474);
   U763 : EOI port map( A => n301, B => n507, Z => n1044);
   U764 : EOI port map( A => n850, B => n633, Z => n507);
   U765 : ENI port map( A => n1073, B => n4735, Z => n475);
   U767 : ENI port map( A => n851, B => n1075, Z => n766);
   U768 : EOI port map( A => n975, B => n339, Z => n1075);
   U769 : ENI port map( A => n898, B => n4736, Z => n339);
   U770 : EOI port map( A => n303, B => n1076, Z => n1071);
   U771 : EOI port map( A => n400, B => n271, Z => n1076);
   U772 : EOI port map( A => n4550, B => n4799, Z => n271);
   U773 : EOI port map( A => n1079, B => n1080, Z => n1069);
   U774 : EOI port map( A => n481, B => n480, Z => n1080);
   U775 : ENI port map( A => n219, B => n1049, Z => n480);
   U776 : EOI port map( A => n307, B => n511, Z => n1049);
   U777 : EOI port map( A => n861, B => n642, Z => n511);
   U778 : ENI port map( A => n1081, B => n4739, Z => n481);
   U780 : ENI port map( A => n862, B => n1083, Z => n773);
   U781 : EOI port map( A => n992, B => n347, Z => n1083);
   U782 : ENI port map( A => n906, B => n4740, Z => n347);
   U783 : EOI port map( A => n309, B => n1084, Z => n1079);
   U784 : EOI port map( A => n406, B => n277, Z => n1084);
   U785 : EOI port map( A => n4449, B => n4799, Z => n277);
   U786 : EOI port map( A => n1086, B => n1087, Z => n1067);
   U787 : EOI port map( A => n313, B => n1088, Z => n1087);
   U788 : EOI port map( A => n412, B => n281, Z => n1088);
   U789 : EOI port map( A => n4446, B => n4799, Z => n281);
   U790 : EOI port map( A => n487, B => n488, Z => n1086);
   U791 : ENI port map( A => n1090, B => n4737, Z => n488);
   U793 : ENI port map( A => n867, B => n1092, Z => n781);
   U794 : EOI port map( A => n983, B => n353, Z => n1092);
   U795 : ENI port map( A => n917, B => n4738, Z => n353);
   U796 : EOI port map( A => n226, B => n1056, Z => n487);
   U797 : EOI port map( A => n316, B => n516, Z => n1056);
   U798 : EOI port map( A => n866, B => n647, Z => n516);
   U800 : EOI port map( A => n1095, B => n1096, Z => n1094);
   U801 : EOI port map( A => n289, B => n1097, Z => n1096);
   U802 : EOI port map( A => n420, B => n321, Z => n1097);
   U803 : EOI port map( A => n4566, B => n4799, Z => n289);
   U804 : EOI port map( A => n495, B => n496, Z => n1095);
   U805 : ENI port map( A => n790, B => n4764, Z => n496);
   U807 : ENI port map( A => n878, B => n1101, Z => n790);
   U808 : EOI port map( A => n4751, B => n360, Z => n1101);
   U809 : EOI port map( A => n928, B => n1102, Z => n360);
   U810 : ENI port map( A => n233, B => n1063, Z => n495);
   U811 : EOI port map( A => n324, B => n522, Z => n1063);
   U812 : EOI port map( A => n880, B => n658, Z => n522);
   U813 : EOI port map( A => n4660, B => v_DATA_COLUMN_13_port, Z => n1093);
   U817 : EOI port map( A => n1110, B => n1111, Z => n1109);
   U818 : EOI port map( A => n301, B => n508, Z => n1111);
   U819 : ENI port map( A => n1112, B => n765, Z => n508);
   U820 : ENI port map( A => n1113, B => n1114, Z => n765);
   U821 : EOI port map( A => n1115, B => n1116, Z => n1114);
   U822 : EOI port map( A => n634, B => n848, Z => n1116);
   U823 : EOI port map( A => n437, B => n4743, Z => n848);
   U825 : EOI port map( A => n3932, B => n4787, Z => n437);
   U826 : ENI port map( A => n1119, B => n847, Z => n1113);
   U827 : ENI port map( A => n121, B => n676, Z => n847);
   U828 : ENI port map( A => n1073, B => n711, Z => n1112);
   U829 : ENI port map( A => n476, B => n303, Z => n711);
   U830 : EOI port map( A => n3919, B => n4664, Z => n303);
   U831 : EOI port map( A => n4547, B => n4760, Z => n476);
   U832 : ENI port map( A => n534, B => n1122, Z => n1073);
   U833 : EOI port map( A => n154, B => n336, Z => n1122);
   U834 : EOI port map( A => n673, B => n402, Z => n154);
   U835 : EOI port map( A => n900, B => n633, Z => n534);
   U836 : ENI port map( A => n4800, B => n160, Z => n301);
   U838 : ENI port map( A => n4444, B => n4659, Z => n338);
   U839 : EOI port map( A => n477, B => n768, Z => n1110);
   U840 : EOI port map( A => n536, B => n161, Z => n768);
   U841 : EOI port map( A => n3911, B => n4669, Z => n477);
   U842 : EOI port map( A => n1124, B => n1125, Z => n1108);
   U843 : EOI port map( A => n307, B => n512, Z => n1125);
   U844 : ENI port map( A => n1126, B => n772, Z => n512);
   U845 : ENI port map( A => n1127, B => n1128, Z => n772);
   U846 : EOI port map( A => n1129, B => n1130, Z => n1128);
   U847 : EOI port map( A => n643, B => n859, Z => n1130);
   U848 : EOI port map( A => n445, B => n4745, Z => n859);
   U850 : EOI port map( A => n3868, B => n4787, Z => n445);
   U851 : ENI port map( A => n1132, B => n858, Z => n1127);
   U852 : ENI port map( A => n127, B => n683, Z => n858);
   U853 : ENI port map( A => n1081, B => n716, Z => n1126);
   U854 : ENI port map( A => n482, B => n309, Z => n716);
   U855 : EOI port map( A => n3855, B => n4664, Z => n309);
   U856 : EOI port map( A => n4447, B => n4760, Z => n482);
   U857 : ENI port map( A => n541, B => n1134, Z => n1081);
   U858 : EOI port map( A => n184, B => n344, Z => n1134);
   U859 : EOI port map( A => n680, B => n408, Z => n184);
   U860 : EOI port map( A => n908, B => n642, Z => n541);
   U861 : ENI port map( A => n4801, B => n181, Z => n307);
   U863 : ENI port map( A => n4448, B => n4659, Z => n346);
   U864 : EOI port map( A => n483, B => n775, Z => n1124);
   U865 : EOI port map( A => n543, B => n182, Z => n775);
   U866 : EOI port map( A => n3847, B => n4669, Z => n483);
   U867 : EOI port map( A => n1136, B => n1137, Z => n1106);
   U868 : EOI port map( A => n486, B => n778, Z => n1137);
   U869 : EOI port map( A => n548, B => n175, Z => n778);
   U870 : EOI port map( A => n3879, B => n4669, Z => n486);
   U871 : EOI port map( A => n515, B => n316, Z => n1136);
   U872 : ENI port map( A => n4802, B => n174, Z => n316);
   U874 : ENI port map( A => n4455, B => n4659, Z => n352);
   U875 : EOI port map( A => n1139, B => n780, Z => n515);
   U876 : ENI port map( A => n1140, B => n1141, Z => n780);
   U877 : EOI port map( A => n1142, B => n1143, Z => n1141);
   U878 : EOI port map( A => n648, B => n869, Z => n1143);
   U879 : EOI port map( A => n451, B => n4744, Z => n869);
   U881 : EOI port map( A => n3900, B => n4787, Z => n451);
   U882 : ENI port map( A => n1145, B => n868, Z => n1140);
   U883 : ENI port map( A => n131, B => n687, Z => n868);
   U884 : EOI port map( A => n1090, B => n4758, Z => n1139);
   U886 : ENI port map( A => n489, B => n313, Z => n722);
   U887 : EOI port map( A => n3887, B => n4664, Z => n313);
   U888 : EOI port map( A => n4563, B => n4760, Z => n489);
   U889 : ENI port map( A => n546, B => n1147, Z => n1090);
   U890 : EOI port map( A => n168, B => n350, Z => n1147);
   U891 : EOI port map( A => n1054, B => n414, Z => n168);
   U892 : EOI port map( A => n912, B => n647, Z => n546);
   U894 : EOI port map( A => n1150, B => n1151, Z => n1149);
   U895 : EOI port map( A => n494, B => n787, Z => n1151);
   U896 : EOI port map( A => n557, B => n203_port, Z => n787);
   U897 : EOI port map( A => n3815, B => n4669, Z => n494);
   U898 : EOI port map( A => n521, B => n324, Z => n1150);
   U899 : ENI port map( A => n4803, B => n204, Z => n324);
   U901 : ENI port map( A => n4401, B => n4659, Z => n362);
   U902 : EOI port map( A => n1153, B => n789, Z => n521);
   U903 : ENI port map( A => n1154, B => n1155, Z => n789);
   U904 : EOI port map( A => n882, B => n1156, Z => n1155);
   U905 : EOI port map( A => n659, B => n1157, Z => n1156);
   U906 : ENI port map( A => n461, B => n4752, Z => n882);
   U907 : EOI port map( A => n4556, B => n4787, Z => n461);
   U908 : EOI port map( A => n1160, B => n881, Z => n1154);
   U909 : EOI port map( A => n143, B => n696, Z => n881);
   U910 : EOI port map( A => n1100, B => n4759, Z => n1153);
   U912 : ENI port map( A => n497, B => n321, Z => n729);
   U913 : EOI port map( A => n3823, B => n4664, Z => n321);
   U914 : EOI port map( A => n4557, B => n4760, Z => n497);
   U915 : ENI port map( A => n558, B => n1162, Z => n1100);
   U916 : EOI port map( A => n201_port, B => n363, Z => n1162);
   U917 : EOI port map( A => n1061, B => n422, Z => n201_port);
   U918 : EOI port map( A => n922, B => n658, Z => n558);
   U919 : EOI port map( A => v_KEY_COLUMN_12_port, B => v_DATA_COLUMN_12_port, 
                           Z => n1148);
   U923 : EOI port map( A => n1170, B => n1171, Z => n1169);
   U924 : EOI port map( A => n335, B => n533, Z => n1171);
   U925 : ENI port map( A => n1119, B => n1115, Z => n533);
   U926 : EOI port map( A => n435, B => n4795, Z => n1115);
   U928 : EOI port map( A => n806, B => n4766, Z => n1119);
   U929 : EOI port map( A => n4560, B => n4780, Z => n806);
   U930 : ENI port map( A => n1175, B => n844, Z => n335);
   U931 : ENI port map( A => n1176, B => n1177, Z => n844);
   U932 : EOI port map( A => n634, B => n1178, Z => n1177);
   U933 : EOI port map( A => n120, B => n899, Z => n1178);
   U934 : EOI port map( A => n158, B => n161, Z => n899);
   U935 : ENI port map( A => n604, B => n804, Z => n1176);
   U936 : EOI port map( A => n4805, B => n4736, Z => n804);
   U938 : ENI port map( A => n4545, B => v_KEY_COLUMN_0_port, Z => n157);
   U939 : EOI port map( A => n4775, B => n536, Z => n1175);
   U940 : EOI port map( A => n4540, B => n4788, Z => n536);
   U942 : ENI port map( A => n4451, B => n4668, Z => n850);
   U943 : EOI port map( A => n336, B => n1185, Z => n1170);
   U944 : EOI port map( A => n846, B => n851, Z => n1185);
   U945 : EOI port map( A => n574, B => n161, Z => n851);
   U946 : EOI port map( A => n4546, B => n4761, Z => n846);
   U947 : EOI port map( A => n438, B => n160, Z => n336);
   U948 : ENI port map( A => n4532, B => n4658, Z => n438);
   U949 : EOI port map( A => n1189, B => n1190, Z => n1168);
   U950 : EOI port map( A => n343, B => n540, Z => n1190);
   U951 : ENI port map( A => n1132, B => n1129, Z => n540);
   U952 : EOI port map( A => n443, B => n4796, Z => n1129);
   U954 : EOI port map( A => n814, B => n4767, Z => n1132);
   U955 : EOI port map( A => n4442, B => n4780, Z => n814);
   U956 : ENI port map( A => n1193, B => n855, Z => n343);
   U957 : ENI port map( A => n1194, B => n1195, Z => n855);
   U958 : EOI port map( A => n643, B => n1196, Z => n1195);
   U959 : EOI port map( A => n126, B => n907, Z => n1196);
   U960 : EOI port map( A => n4793, B => n4783, Z => n907);
   U962 : ENI port map( A => n608, B => n812, Z => n1194);
   U963 : EOI port map( A => n185, B => n639, Z => n812);
   U964 : EOI port map( A => n4553, B => n4804, Z => n185);
   U965 : EOI port map( A => n4776, B => n543, Z => n1193);
   U966 : EOI port map( A => n4536, B => n4788, Z => n543);
   U968 : ENI port map( A => n4443, B => n4668, Z => n861);
   U969 : EOI port map( A => n344, B => n1203, Z => n1189);
   U970 : EOI port map( A => n857, B => n862, Z => n1203);
   U971 : EOI port map( A => n580, B => n182, Z => n862);
   U972 : EOI port map( A => n4554, B => n4761, Z => n857);
   U973 : EOI port map( A => n446, B => n181, Z => n344);
   U974 : ENI port map( A => n4533, B => n4658, Z => n446);
   U975 : EOI port map( A => n1206, B => n1207, Z => n1166);
   U976 : EOI port map( A => n350, B => n1208, Z => n1207);
   U977 : EOI port map( A => n873, B => n867, Z => n1208);
   U978 : EOI port map( A => n584, B => n175, Z => n867);
   U979 : EOI port map( A => n4562, B => n4761, Z => n873);
   U980 : EOI port map( A => n452, B => n174, Z => n350);
   U981 : ENI port map( A => n4432, B => n4658, Z => n452);
   U982 : EOI port map( A => n549, B => n354, Z => n1206);
   U983 : ENI port map( A => n1211, B => n871, Z => n354);
   U984 : ENI port map( A => n1212, B => n1213, Z => n871);
   U985 : EOI port map( A => n648, B => n1214, Z => n1213);
   U986 : EOI port map( A => n130, B => n914, Z => n1214);
   U987 : EOI port map( A => n172, B => n175, Z => n914);
   U988 : EOI port map( A => n954, B => n821, Z => n1212);
   U989 : EOI port map( A => n4806, B => n4738, Z => n821);
   U991 : ENI port map( A => n4561, B => v_KEY_COLUMN_0_port, Z => n171);
   U992 : EOI port map( A => n4777, B => n548, Z => n1211);
   U993 : EOI port map( A => n4552, B => n4788, Z => n548);
   U995 : ENI port map( A => n4453, B => n4668, Z => n866);
   U996 : EOI port map( A => n1145, B => n1142, Z => n549);
   U997 : EOI port map( A => n449, B => n414, Z => n1142);
   U998 : EOI port map( A => n817, B => n4768, Z => n1145);
   U999 : EOI port map( A => n4543, B => n4780, Z => n817);
   U1001 : EOI port map( A => n1223, B => n1224, Z => n1222);
   U1002 : EOI port map( A => n878, B => n1225, Z => n1224);
   U1003 : EOI port map( A => n886, B => n363, Z => n1225);
   U1004 : EOI port map( A => n462, B => n204, Z => n363);
   U1005 : EOI port map( A => n4430, B => n4390, Z => n462);
   U1006 : EOI port map( A => n4538, B => n4761, Z => n886);
   U1007 : EOI port map( A => n592, B => n203_port, Z => n878);
   U1008 : EOI port map( A => n561, B => n365, Z => n1223);
   U1009 : ENI port map( A => n1229, B => n884, Z => n365);
   U1010 : ENI port map( A => n1230, B => n1231, Z => n884);
   U1011 : EOI port map( A => n659, B => n1232, Z => n1231);
   U1012 : EOI port map( A => n141, B => n924, Z => n1232);
   U1013 : EOI port map( A => n189, B => n203_port, Z => n924);
   U1014 : EOI port map( A => n964, B => n832, Z => n1230);
   U1015 : EOI port map( A => n4807, B => n4742, Z => n832);
   U1017 : ENI port map( A => n4555, B => v_KEY_COLUMN_0_port, Z => n656);
   U1018 : EOI port map( A => n4778, B => n557, Z => n1229);
   U1019 : EOI port map( A => n4531, B => n4788, Z => n557);
   U1021 : ENI port map( A => n4436, B => n4668, Z => n880);
   U1022 : EOI port map( A => n1160, B => n1157, Z => n561);
   U1023 : EOI port map( A => n459, B => n422, Z => n1157);
   U1024 : EOI port map( A => n4781, B => n1061, Z => n1160);
   U1026 : ENI port map( A => n4558, B => v_KEY_COLUMN_25_port, Z => n827);
   U1027 : EOI port map( A => n4659, B => v_DATA_COLUMN_11_port, Z => n1221);
   U1031 : EOI port map( A => n1246, B => n1247, Z => n1245);
   U1032 : EOI port map( A => n571, B => n803, Z => n1247);
   U1033 : EOI port map( A => n435, B => n4790, Z => n803);
   U1035 : ENI port map( A => n4568, B => n4663, Z => n121);
   U1036 : EOI port map( A => n3924, B => n4725, Z => n435);
   U1037 : EOI port map( A => n604, B => n120, Z => n571);
   U1038 : EOI port map( A => n977, B => n160, Z => n120);
   U1039 : ENI port map( A => n1251, B => n633, Z => n604);
   U1040 : EOI port map( A => n898, B => n434, Z => n1246);
   U1041 : ENI port map( A => n1252, B => n897, Z => n434);
   U1042 : EOI port map( A => n801, B => n118, Z => n897);
   U1043 : ENI port map( A => n1253, B => n1254, Z => n118);
   U1044 : EOI port map( A => n160, B => n402, Z => n1254);
   U1045 : ENI port map( A => n4431, B => n4661, Z => n402);
   U1046 : EOI port map( A => n4766, B => n633, Z => n1253);
   U1047 : EOI port map( A => n3914, B => n4671, Z => n633);
   U1049 : ENI port map( A => n4438, B => n4670, Z => n673);
   U1050 : ENI port map( A => n1257, B => n975, Z => n801);
   U1051 : EOI port map( A => n4736, B => n161, Z => n1257);
   U1052 : ENI port map( A => n4525, B => n4666, Z => n161);
   U1054 : ENI port map( A => n900, B => n574, Z => n1252);
   U1055 : EOI port map( A => n4539, B => n4789, Z => n574);
   U1056 : EOI port map( A => n4541, B => n4779, Z => n900);
   U1057 : EOI port map( A => n4517, B => n4771, Z => n898);
   U1059 : EOI port map( A => n577, B => n811, Z => n1266);
   U1060 : EOI port map( A => n443, B => n4791, Z => n811);
   U1062 : ENI port map( A => n4567, B => n4663, Z => n127);
   U1063 : EOI port map( A => n3860, B => n4725, Z => n443);
   U1064 : EOI port map( A => n608, B => n126, Z => n577);
   U1065 : EOI port map( A => n990, B => n181, Z => n126);
   U1066 : ENI port map( A => n1269, B => n642, Z => n608);
   U1067 : EOI port map( A => n906, B => n442, Z => n1265);
   U1068 : ENI port map( A => n1270, B => n905, Z => n442);
   U1069 : EOI port map( A => n809, B => n124, Z => n905);
   U1070 : ENI port map( A => n1271, B => n1272, Z => n124);
   U1071 : EOI port map( A => n181, B => n408, Z => n1272);
   U1072 : ENI port map( A => n4434, B => n4661, Z => n408);
   U1073 : EOI port map( A => n4767, B => n642, Z => n1271);
   U1074 : EOI port map( A => n3850, B => n4671, Z => n642);
   U1076 : ENI port map( A => n4428, B => n4670, Z => n680);
   U1077 : ENI port map( A => n1275, B => n992, Z => n809);
   U1078 : EOI port map( A => n4740, B => n182, Z => n1275);
   U1079 : ENI port map( A => n4522, B => n4666, Z => n182);
   U1081 : ENI port map( A => n908, B => n580, Z => n1270);
   U1082 : EOI port map( A => n4535, B => n4789, Z => n580);
   U1083 : EOI port map( A => n4528, B => n4779, Z => n908);
   U1084 : EOI port map( A => n4421, B => n4771, Z => n906);
   U1086 : EOI port map( A => n1280, B => n1281, Z => n1242);
   U1087 : EOI port map( A => n917, B => n453, Z => n1281);
   U1088 : ENI port map( A => n1282, B => n916, Z => n453);
   U1089 : EOI port map( A => n818, B => n133, Z => n916);
   U1090 : ENI port map( A => n1283, B => n1284, Z => n133);
   U1091 : EOI port map( A => n174, B => n414, Z => n1284);
   U1092 : ENI port map( A => n4433, B => n4661, Z => n414);
   U1093 : EOI port map( A => n4768, B => n647, Z => n1283);
   U1095 : ENI port map( A => n4427, B => n4670, Z => n1054);
   U1096 : ENI port map( A => n1287, B => n983, Z => n818);
   U1097 : EOI port map( A => n4738, B => n175, Z => n1287);
   U1098 : ENI port map( A => n4420, B => n4666, Z => n175);
   U1100 : ENI port map( A => n912, B => n584, Z => n1282);
   U1101 : EOI port map( A => n4551, B => n4789, Z => n584);
   U1102 : EOI port map( A => n4544, B => n4779, Z => n912);
   U1103 : EOI port map( A => n4542, B => n4771, Z => n917);
   U1104 : ENI port map( A => n820, B => n586, Z => n1280);
   U1105 : EOI port map( A => n4762, B => n130, Z => n586);
   U1106 : EOI port map( A => n985, B => n174, Z => n130);
   U1108 : EOI port map( A => n1293, B => n647, Z => n954);
   U1109 : EOI port map( A => n3882, B => n4671, Z => n647);
   U1110 : ENI port map( A => n4726, B => n131, Z => n820);
   U1111 : ENI port map( A => n4570, B => n4663, Z => n131);
   U1113 : ENI port map( A => n4445, B => v_KEY_COLUMN_9_port, Z => n449);
   U1115 : EOI port map( A => n1299, B => n1300, Z => n1298);
   U1116 : EOI port map( A => n928, B => n464, Z => n1300);
   U1117 : ENI port map( A => n1301, B => n926, Z => n464);
   U1118 : EOI port map( A => n828, B => n140, Z => n926);
   U1119 : ENI port map( A => n1302, B => n1303, Z => n140);
   U1120 : EOI port map( A => n422, B => n658, Z => n1303);
   U1121 : ENI port map( A => n4398, B => n4661, Z => n422);
   U1122 : EOI port map( A => n204, B => n4769, Z => n1302);
   U1124 : ENI port map( A => n4437, B => n4670, Z => n1061);
   U1125 : ENI port map( A => n1306, B => n1307, Z => n828);
   U1126 : EOI port map( A => n203_port, B => n696, Z => n1307);
   U1127 : EOI port map( A => n4518, B => n4387, Z => n203_port);
   U1128 : EOI port map( A => n4742, B => n231, Z => n1306);
   U1129 : ENI port map( A => n592, B => n922, Z => n1301);
   U1130 : EOI port map( A => n4559, B => n4779, Z => n922);
   U1131 : EOI port map( A => n4549, B => n4789, Z => n592);
   U1132 : ENI port map( A => n4537, B => v_KEY_COLUMN_2_port, Z => n928);
   U1133 : EOI port map( A => n831, B => n594, Z => n1299);
   U1134 : EOI port map( A => n4763, B => n141, Z => n594);
   U1135 : EOI port map( A => n995, B => n204, Z => n141);
   U1137 : EOI port map( A => n1313, B => n658, Z => n964);
   U1138 : EOI port map( A => n3818, B => n4671, Z => n658);
   U1139 : EOI port map( A => n4728, B => n143, Z => n831);
   U1140 : EOI port map( A => n4548, B => n4403, Z => n143);
   U1142 : ENI port map( A => n4429, B => v_KEY_COLUMN_9_port, Z => n459);
   U1143 : EOI port map( A => n4658, B => v_DATA_COLUMN_10_port, Z => n1297);
   U1145 : AO1P port map( A => n1321, B => n4386, C => n1322, D => n1323, Z => 
                           n1320);
   U1146 : NR2I port map( A => n4383, B => n1324, Z => n1323);
   U1147 : EOI port map( A => n1325, B => n1326, Z => n1324);
   U1148 : EOI port map( A => n671, B => n629, Z => n1326);
   U1149 : EOI port map( A => n158, B => n977, Z => n629);
   U1150 : EOI port map( A => n4519, B => n4732, Z => n977);
   U1151 : EOI port map( A => n4523, B => n4792, Z => n158);
   U1152 : EOI port map( A => n631, B => n160, Z => n671);
   U1153 : EOI port map( A => n3930, B => n4662, Z => n160);
   U1154 : ENI port map( A => n4417, B => n4657, Z => n631);
   U1155 : EOI port map( A => n156, B => n975, Z => n1325);
   U1156 : EOI port map( A => n676, B => n216, Z => n975);
   U1157 : ENI port map( A => n4416, B => n4656, Z => n216);
   U1158 : EOI port map( A => n3921, B => n4665, Z => n676);
   U1159 : ENI port map( A => n1251, B => n634, Z => n156);
   U1160 : ENI port map( A => n214, B => n376, Z => n634);
   U1161 : EOI port map( A => n400, B => n243, Z => n376);
   U1162 : EOI port map( A => n3928, B => n4660, Z => n243);
   U1163 : EOI port map( A => n4510, B => n4773, Z => n400);
   U1164 : ENI port map( A => n270, B => n403, Z => n214);
   U1165 : EOI port map( A => n3936, B => n4655, Z => n403);
   U1166 : EOI port map( A => n4524, B => n4785, Z => n270);
   U1167 : EOI port map( A => n4456, B => n4667, Z => n1251);
   U1170 : EOI port map( A => n1341, B => n1342, Z => n1340);
   U1171 : EOI port map( A => n689, B => n650, Z => n1342);
   U1172 : EOI port map( A => n172, B => n985, Z => n650);
   U1173 : EOI port map( A => n4419, B => n4732, Z => n985);
   U1174 : EOI port map( A => n4520, B => n4792, Z => n172);
   U1175 : EOI port map( A => n1289, B => n174, Z => n689);
   U1176 : EOI port map( A => n3898, B => n4662, Z => n174);
   U1177 : ENI port map( A => n4439, B => n4657, Z => n1289);
   U1178 : EOI port map( A => n170, B => n983, Z => n1341);
   U1179 : EOI port map( A => n687, B => n224, Z => n983);
   U1180 : ENI port map( A => n4425, B => n4656, Z => n224);
   U1181 : EOI port map( A => n3889, B => n4665, Z => n687);
   U1182 : ENI port map( A => n1293, B => n648, Z => n170);
   U1183 : EOI port map( A => n4753, B => n384, Z => n648);
   U1184 : EOI port map( A => n412, B => n251, Z => n384);
   U1185 : EOI port map( A => n3896, B => n4660, Z => n251);
   U1186 : EOI port map( A => n4507, B => n4773, Z => n412);
   U1188 : ENI port map( A => n280, B => n415, Z => n226);
   U1189 : EOI port map( A => n3904, B => n4655, Z => n415);
   U1190 : EOI port map( A => n4415, B => n4785, Z => n280);
   U1191 : EOI port map( A => n4440, B => n4667, Z => n1293);
   U1196 : EOI port map( A => v_DATA_COLUMN_0_port, B => n4804, Z => n1339);
   U1199 : EOI port map( A => n1355, B => n1356, Z => n1321);
   U1200 : EOI port map( A => n186, B => n992, Z => n1356);
   U1201 : EOI port map( A => n683, B => n221, Z => n992);
   U1202 : ENI port map( A => n4397, B => n4656, Z => n221);
   U1203 : EOI port map( A => n3857, B => n4665, Z => n683);
   U1204 : ENI port map( A => n1269, B => n643, Z => n186);
   U1205 : ENI port map( A => n219, B => n380, Z => n643);
   U1206 : EOI port map( A => n406, B => n247, Z => n380);
   U1207 : EOI port map( A => n3864, B => n4660, Z => n247);
   U1208 : EOI port map( A => n4413, B => n4773, Z => n406);
   U1209 : ENI port map( A => n276, B => n409, Z => n219);
   U1210 : EOI port map( A => n3872, B => n4655, Z => n409);
   U1211 : EOI port map( A => n4521, B => n4785, Z => n276);
   U1212 : EOI port map( A => n4454, B => n4667, Z => n1269);
   U1213 : EOI port map( A => n640, B => n678, Z => n1355);
   U1214 : EOI port map( A => n639, B => n181, Z => n678);
   U1215 : EOI port map( A => n3866, B => n4662, Z => n181);
   U1216 : ENI port map( A => n4422, B => n4657, Z => n639);
   U1217 : EOI port map( A => n4793, B => n990, Z => n640);
   U1218 : EOI port map( A => n4423, B => n4732, Z => n990);
   U1220 : ENI port map( A => n4534, B => v_KEY_COLUMN_16_port, Z => n179);
   U1228 : ENI port map( A => n4794, B => n995, Z => n661);
   U1229 : ENI port map( A => n4529, B => v_KEY_COLUMN_8_port, Z => n995);
   U1231 : ENI port map( A => n4530, B => v_KEY_COLUMN_16_port, Z => n189);
   U1234 : ND2I port map( A => n4382, B => n4756, Z => n199_port);
   U1237 : EOI port map( A => n4752, B => n696, Z => n1371);
   U1239 : ENI port map( A => n4424, B => n4656, Z => n231);
   U1240 : ND2I port map( A => n1376, B => n4382, Z => n197);
   U1245 : EOI port map( A => n1313, B => n659, Z => n1376);
   U1246 : EOI port map( A => n390, B => n233, Z => n659);
   U1247 : EOI port map( A => n4786, B => n4757, Z => n233);
   U1248 : EOI port map( A => n258, B => n420, Z => n390);
   U1249 : EOI port map( A => n3816, B => v_KEY_COLUMN_29_port, Z => n420);
   U1250 : EOI port map( A => n4414, B => n4385, Z => n258);
   U1251 : EOI port map( A => n4450, B => n4667, Z => n1313);
   U1252 : EOI port map( A => n4742, B => n204, Z => n1364);
   U1253 : EOI port map( A => n4418, B => n4388, Z => n204);
   U1255 : ENI port map( A => n4435, B => n4657, Z => n1102);
   U1261 : ND2I port map( A => N203, B => n1392, Z => n1394);
   U1263 : ND2I port map( A => N202, B => n1392, Z => n1395);
   U1265 : ND2I port map( A => N201, B => n1392, Z => n1396);
   U1269 : ND2I port map( A => N199, B => n1392, Z => n1399);
   U1271 : ND2I port map( A => n4620, B => n1392, Z => n1400);
   U1308 : ND2I port map( A => n1425, B => v_CNT4_0_port, Z => n1415);
   U1343 : ND2I port map( A => n1444, B => n4395, Z => n1408);
   U1345 : ND2I port map( A => n4589, B => CE_I, Z => n1445);
   U1347 : ND2I port map( A => v_CNT4_0_port, B => n1444, Z => n1404);
   U1348 : NR2I port map( A => n4840, B => v_CNT4_1_port, Z => n1444);
   U1350 : ND2I port map( A => CE_I, B => n4395, Z => n1447);
   U1566 : ND2I port map( A => n1471, B => n4463, Z => n1476);
   U1572 : NR2I port map( A => n4845, B => n4853, Z => n1477);
   U1575 : ND2I port map( A => n4850, B => n1482, Z => n1480);
   U1583 : AO1P port map( A => n3946, B => n4854, C => n1487, D => n1467, Z => 
                           n4300);
   U1584 : NR2I port map( A => n4854, B => n3946, Z => n1467);
   U1586 : ND2I port map( A => n3956, B => VALID_DATA_I, Z => n1398);
   U1588 : NR2I port map( A => n4713, B => n3947, Z => n1465);
   U1589 : ND2I port map( A => n1489, B => n1490, Z => n4291);
   U1591 : NR2I port map( A => v_CALCULATION_CNTR_3_port, B => 
                           v_CALCULATION_CNTR_2_port, Z => n1492);
   U1596 : ND2I port map( A => n1494, B => n1495, Z => n4292);
   U1600 : ND2I port map( A => n3940, B => CE_I, Z => n103);
   U1616 : ND2I port map( A => n1528, B => n4599, Z => n1524);
   U1620 : ND2I port map( A => n1534, B => n4434, Z => n1531);
   U1624 : ND2I port map( A => n1539, B => n4598, Z => n1536);
   U1628 : ND2I port map( A => n1543, B => n4449, Z => n1541);
   U1632 : ND2I port map( A => n1548, B => n4448, Z => n1545);
   U1636 : ND2I port map( A => n1552, B => n4533, Z => n1550);
   U1640 : ND2I port map( A => n1557, B => n4597, Z => n1554);
   U1644 : ND2I port map( A => n1561, B => n4423, Z => n1559);
   U1646 : ND2I port map( A => n1529, B => n1527, Z => n1523);
   U1647 : ND2I port map( A => n1527, B => n1562, Z => n1529);
   U1650 : ND2I port map( A => n1568, B => n4422, Z => n1565);
   U1654 : ND2I port map( A => n1574, B => n4397, Z => n1571);
   U1658 : ND2I port map( A => n1580, B => n4596, Z => n1576);
   U1662 : ND2I port map( A => n1584, B => n4447, Z => n1582);
   U1666 : ND2I port map( A => n1588, B => n4554, Z => n1586);
   U1670 : ND2I port map( A => n1592, B => n4421, Z => n1590);
   U1674 : ND2I port map( A => n1597, B => n4595, Z => n1594);
   U1678 : ND2I port map( A => n1601, B => n4553, Z => n1599);
   U1680 : ND2I port map( A => n1569, B => n1527, Z => n1564);
   U1681 : ND2I port map( A => n1527, B => n1602, Z => n1569);
   U1684 : ND2I port map( A => n1610, B => n4591, Z => n1605);
   U1688 : ND2I port map( A => n1616, B => n4427, Z => n1613);
   U1692 : ND2I port map( A => n1620, B => n4507, Z => n1618);
   U1696 : ND2I port map( A => n1626, B => n4590, Z => n1622);
   U1700 : ND2I port map( A => n1631, B => n4453, Z => n1628);
   U1704 : ND2I port map( A => n1635, B => n4544, Z => n1633);
   U1708 : ND2I port map( A => n1639, B => n4543, Z => n1637);
   U1712 : ND2I port map( A => n1644, B => n4440, Z => n1641);
   U1714 : ND2I port map( A => n1611, B => n1609, Z => n1604);
   U1715 : ND2I port map( A => n1609, B => n1602, Z => n1611);
   U1718 : ND2I port map( A => n1649, B => n4420, Z => n1647);
   U1722 : ND2I port map( A => n1656, B => n4583, Z => n1652);
   U1726 : ND2I port map( A => n1660, B => n4415, Z => n1658);
   U1730 : ND2I port map( A => n1666, B => n4582, Z => n1662);
   U1734 : ND2I port map( A => n1670, B => n4552, Z => n1668);
   U1737 : ND2I port map( A => n1674, B => n4551, Z => n1673);
   U1743 : ND2I port map( A => n1685, B => n1686, Z => n1684);
   U1748 : ND2I port map( A => n1697, B => n4570, Z => n1695);
   U1751 : ND2I port map( A => n1701, B => n4520, Z => n1700);
   U1754 : ND2I port map( A => n1650, B => n1609, Z => n1646);
   U1755 : ND2I port map( A => n1609, B => n1702, Z => n1650);
   U1768 : ND2I port map( A => n1730, B => n4581, Z => n1727);
   U1772 : ND2I port map( A => n1734, B => n4433, Z => n1732);
   U1776 : ND2I port map( A => n1738, B => n4580, Z => n1735);
   U1780 : ND2I port map( A => n1741, B => n4446, Z => n1739);
   U1784 : ND2I port map( A => n1744, B => n4455, Z => n1742);
   U1788 : ND2I port map( A => n1747, B => n4432, Z => n1745);
   U1792 : ND2I port map( A => n1750, B => n4445, Z => n1748);
   U1796 : ND2I port map( A => n1753, B => n4419, Z => n1751);
   U1798 : ND2I port map( A => n1731, B => n1609, Z => n1726);
   U1799 : ND2I port map( A => n1609, B => n1754, Z => n1731);
   U1802 : ND2I port map( A => n1758, B => n4439, Z => n1756);
   U1807 : ND2I port map( A => n1762, B => n4425, Z => n1760);
   U1812 : ND2I port map( A => n1766, B => n4618, Z => n1763);
   U1817 : ND2I port map( A => n1769, B => n4563, Z => n1767);
   U1822 : ND2I port map( A => n1772, B => n4562, Z => n1770);
   U1827 : ND2I port map( A => n1775, B => n4542, Z => n1773);
   U1832 : ND2I port map( A => n1779, B => n4617, Z => n1776);
   U1837 : ND2I port map( A => n1782, B => n4561, Z => n1780);
   U1840 : ND2I port map( A => n1759, B => n1609, Z => n1755);
   U1841 : ND2I port map( A => n1609, B => n1562, Z => n1759);
   U1844 : ND2I port map( A => n1787, B => n4616, Z => n1784);
   U1849 : ND2I port map( A => n1791, B => n4438, Z => n1789);
   U1854 : ND2I port map( A => n1794, B => n4510, Z => n1792);
   U1859 : ND2I port map( A => n1798, B => n4615, Z => n1795);
   U1864 : ND2I port map( A => n1801, B => n4451, Z => n1799);
   U1869 : ND2I port map( A => n1804, B => n4541, Z => n1802);
   U1874 : ND2I port map( A => n1807, B => n4560, Z => n1805);
   U1879 : ND2I port map( A => n1810, B => n4456, Z => n1808);
   U1882 : ND2I port map( A => n1788, B => n4352, Z => n1783);
   U1883 : ND2I port map( A => n4352, B => n1562, Z => n1788);
   U1886 : ND2I port map( A => n1814, B => n4525, Z => n1812);
   U1891 : ND2I port map( A => n1819, B => n4614, Z => n1816);
   U1896 : ND2I port map( A => n1822, B => n4524, Z => n1820);
   U1901 : ND2I port map( A => n1826, B => n4613, Z => n1823);
   U1906 : ND2I port map( A => n1829, B => n4540, Z => n1827);
   U1911 : ND2I port map( A => n1833, B => n4539, Z => n1831);
   U1916 : ND2I port map( A => n1836, B => n4568, Z => n1834);
   U1921 : ND2I port map( A => n1840, B => n4523, Z => n1838);
   U1924 : ND2I port map( A => n1815, B => n4352, Z => n1811);
   U1925 : ND2I port map( A => n4352, B => n1602, Z => n1815);
   U1928 : ND2I port map( A => n1845, B => n4607, Z => n1842);
   U1932 : ND2I port map( A => n1849, B => n4431, Z => n1847);
   U1936 : ND2I port map( A => n1853, B => n4606, Z => n1850);
   U1940 : ND2I port map( A => n1856, B => n4550, Z => n1854);
   U1944 : ND2I port map( A => n1859, B => n4444, Z => n1857);
   U1948 : ND2I port map( A => n1863, B => n4532, Z => n1861);
   U1953 : ND2I port map( A => n4987, B => n5041, Z => n1872);
   U1955 : ND2I port map( A => n5040, B => n4976, Z => n1879);
   U1958 : ND2I port map( A => n1885, B => n4605, Z => n1882);
   U1961 : ND2I port map( A => n1889, B => n4519, Z => n1888);
   U1964 : ND2I port map( A => n1846, B => n4352, Z => n1841);
   U1965 : ND2I port map( A => n4352, B => n1702, Z => n1846);
   U1969 : ND2I port map( A => n1900, B => n1901, Z => n1899);
   U1972 : NR2I port map( A => n1909, B => n1901, Z => n1893);
   U1978 : ND2I port map( A => n1922, B => n4612, Z => n1918);
   U1983 : ND2I port map( A => n1926, B => n4437, Z => n1924);
   U1988 : ND2I port map( A => n1930, B => n4611, Z => n1927);
   U1993 : ND2I port map( A => n1934, B => n4610, Z => n1931);
   U1998 : ND2I port map( A => n1937, B => n4436, Z => n1935);
   U2003 : ND2I port map( A => n1940, B => n4559, Z => n1938);
   U2009 : AO1P port map( A => n4913, B => n1951, C => n1952, D => n1953, Z => 
                           n1948);
   U2010 : NR2I port map( A => n4705, B => n1955, Z => n1953);
   U2014 : ND2I port map( A => n1962, B => n4558, Z => n1960);
   U2019 : ND2I port map( A => n1965, B => n4450, Z => n1963);
   U2022 : ND2I port map( A => n1923, B => n4706, Z => n1917);
   U2023 : ND2I port map( A => n4706, B => n1754, Z => n1923);
   U2026 : AO1P port map( A => n5059, B => n4686, C => n1974, D => n1975, Z => 
                           n1969);
   U2027 : AN2I port map( A => n5061, B => n1977, Z => n1975);
   U2036 : ND2I port map( A => n1994, B => n4518, Z => n1992);
   U2041 : ENI port map( A => n4526, B => n4665, Z => n696);
   U2045 : ENI port map( A => n4514, B => v_KEY_COLUMN_21_port, Z => n288);
   U2048 : ND2I port map( A => n2005, B => n4594, Z => n2002);
   U2052 : ND2I port map( A => n2008, B => n4531, Z => n2006);
   U2056 : ND2I port map( A => n2011, B => n4549, Z => n2009);
   U2060 : ND2I port map( A => n2014, B => n4548, Z => n2012);
   U2064 : ND2I port map( A => n2017, B => n4530, Z => n2015);
   U2066 : ND2I port map( A => n1995, B => n4706, Z => n1991);
   U2067 : ND2I port map( A => n4706, B => n1562, Z => n1995);
   U2072 : ND2I port map( A => n2023, B => n4418, Z => n2021);
   U2076 : ND2I port map( A => n4906, B => n2031, Z => n2029);
   U2078 : ND2I port map( A => n4979, B => n2035, Z => n2033);
   U2085 : ND2I port map( A => n5040, B => n4980, Z => n2052);
   U2089 : ND2I port map( A => n4701, B => n2064, Z => n2057);
   U2091 : AO1P port map( A => n4910, B => n2069, C => n2070, D => n2071, Z => 
                           n2025);
   U2092 : AO1P port map( A => n4702, B => n2072, C => n2073, D => n2074, Z => 
                           n2071);
   U2097 : AO1P port map( A => n2084_port, B => n4701, C => n2085_port, D => 
                           n4962, Z => n2083_port);
   U2100 : AO1P port map( A => n2090, B => n2066, C => n2091, D => n2092, Z => 
                           n2082);
   U2101 : NR2I port map( A => n4955, B => n4361, Z => n2092);
   U2105 : ND2I port map( A => n2096, B => n2097, Z => n2069);
   U2111 : ND2I port map( A => n2103, B => n4398, Z => n2101);
   U2115 : ND2I port map( A => n4506, B => n2109, Z => n2108);
   U2119 : NR2I port map( A => n4971, B => n4966, Z => n2114);
   U2121 : AO1P port map( A => n4971, B => n4701, C => n2118, D => n2119, Z => 
                           n2117);
   U2123 : NR2I port map( A => n4964, B => n4690, Z => n2118);
   U2131 : NR2I port map( A => n4964, B => n4991, Z => n2131);
   U2135 : AO1P port map( A => n4702, B => n2140, C => n2141, D => n2142, Z => 
                           n2139);
   U2136 : NR2I port map( A => n4977, B => n4707, Z => n2142);
   U2138 : AO1P port map( A => n4701, B => n2146, C => n2147, D => n2148, Z => 
                           n2138);
   U2140 : NR2I port map( A => n4965, B => n4984, Z => n2150);
   U2141 : ND2I port map( A => n2153, B => n2154, Z => n2146);
   U2145 : NR2I port map( A => n4980, B => n4977, Z => n2160);
   U2146 : AO1P port map( A => n2113, B => n4379, C => n2163, D => n2164, Z => 
                           n2155);
   U2149 : ND2I port map( A => n2167, B => n2165, Z => n2056);
   U2153 : ND2I port map( A => n2170, B => n4414, Z => n2168);
   U2156 : AO1P port map( A => v_RAM_OUT0_15_port, B => n2173, C => n2174, D =>
                           n2175, Z => n2172);
   U2160 : AO1P port map( A => n4991, B => n4379, C => n2180, D => n2181, Z => 
                           n2174);
   U2166 : ND2I port map( A => n2188, B => n2189, Z => n2187);
   U2169 : NR2I port map( A => n5069, B => n2113, Z => n2129);
   U2170 : AO1P port map( A => n4906, B => n2194, C => n2195, D => n2196, Z => 
                           n2171);
   U2171 : AO1P port map( A => n1916, B => n4360, C => n2197, D => n2198, Z => 
                           n2196);
   U2173 : NR2I port map( A => n4989, B => n4960, Z => n2199);
   U2176 : AO1P port map( A => n4360, B => n2203, C => n2204, D => n2205, Z => 
                           n2202);
   U2178 : NR2I port map( A => n4970, B => n4989, Z => n2206);
   U2179 : AO1P port map( A => n4379, B => n2190, C => n2208, D => n2209, Z => 
                           n2201);
   U2180 : AN2I port map( A => n4360, B => n2210, Z => n2209);
   U2182 : ND2I port map( A => n2213, B => n2214, Z => n2194);
   U2188 : ND2I port map( A => n2219, B => n4566, Z => n2217);
   U2190 : ND2I port map( A => n2220, B => n2221, Z => n1540);
   U2192 : ND2I port map( A => n4910, B => n2225, Z => n2224);
   U2195 : NR2I port map( A => n4976, B => n4955, Z => n2211);
   U2196 : NR2I port map( A => n4983, B => n2095, Z => n2191);
   U2198 : ND2I port map( A => n2232, B => n2233, Z => n2231);
   U2200 : ND2I port map( A => n1914, B => n2226, Z => n2182);
   U2210 : AO1P port map( A => n4506, B => n2250, C => v_RAM_OUT0_9_port, D => 
                           n2251, Z => n2249);
   U2214 : ND2I port map( A => n2256, B => n2257, Z => n2250);
   U2218 : NR2I port map( A => n2061, B => n4963, Z => n2145);
   U2225 : AO1P port map( A => n2264, B => n4379, C => n2265, D => n4702, Z => 
                           n2247);
   U2227 : NR2I port map( A => n4971, B => n4978, Z => n2264);
   U2231 : ND2I port map( A => n2268, B => n4401, Z => n2266);
   U2238 : ND2I port map( A => v_RAM_OUT0_11_port, B => n4391, Z => n2277);
   U2240 : AO1P port map( A => n4968, B => n2281, C => n2282, D => n2241, Z => 
                           n2279);
   U2241 : AN2I port map( A => n2283, B => n4360, Z => n2282);
   U2246 : ND2I port map( A => n4977, B => n2154, Z => n2066);
   U2248 : NR2I port map( A => n4960, B => n4980, Z => n2291);
   U2255 : NR2I port map( A => n2300, B => n2301, Z => n2299);
   U2257 : NR2I port map( A => n4976, B => n2032, Z => n2210);
   U2262 : ND2I port map( A => n2120, B => n2072, Z => n2283);
   U2268 : ND2I port map( A => n2093, B => n1906, Z => n2203);
   U2273 : ND2I port map( A => n2315, B => n4430, Z => n2313);
   U2276 : ND2I port map( A => n4904, B => n1869, Z => n2317);
   U2279 : ND2I port map( A => n2093, B => n2281, Z => n2290);
   U2281 : AO1P port map( A => n4360, B => v_RAM_OUT0_11_port, C => n2324, D =>
                           n2148, Z => n2323);
   U2282 : NR2I port map( A => n2165, B => n4359, Z => n2148);
   U2283 : NR2I port map( A => n4707, B => n2130, Z => n2324);
   U2285 : ND2I port map( A => n2167, B => n2130, Z => n2133);
   U2287 : ND2I port map( A => n2072, B => n2162, Z => n2325);
   U2289 : ND2I port map( A => n4396, B => n4569, Z => n1868);
   U2292 : ND2I port map( A => v_RAM_OUT0_15_port, B => n4569, Z => n2294);
   U2293 : AN2I port map( A => n2329, B => n2330, Z => n1870);
   U2297 : ND2I port map( A => n2212, B => n2162, Z => n2239);
   U2300 : ND2I port map( A => n2281, B => n2212, Z => n2332);
   U2302 : NR2I port map( A => n4987, B => n2113, Z => n2084_port);
   U2306 : AO1P port map( A => n2113, B => n4404, C => n4957, D => n2340, Z => 
                           n2339);
   U2309 : NR2I port map( A => n4691, B => n2342, Z => n2338);
   U2311 : NR2I port map( A => n4994, B => n4991, Z => n2179);
   U2314 : AN2I port map( A => n2344, B => n2226, Z => n2048);
   U2315 : ND2I port map( A => n4960, B => n4702, Z => n2341);
   U2319 : ND2I port map( A => n2120, B => n2347, Z => n2140);
   U2320 : AO1P port map( A => n4988, B => n4379, C => n2349, D => n4968, Z => 
                           n2334);
   U2322 : ND2I port map( A => n4702, B => n2064, Z => n2236);
   U2325 : ND2I port map( A => n4990, B => n4391, Z => n2165);
   U2329 : ND2I port map( A => n2352, B => n4429, Z => n2350);
   U2334 : NR2I port map( A => n2359, B => n2360, Z => n2358);
   U2337 : NR2I port map( A => n4995, B => n4984, Z => n2293);
   U2338 : AO1P port map( A => n4360, B => n2098, C => n2361, D => n2362, Z => 
                           n2357);
   U2342 : NR2I port map( A => n5069, B => n4980, Z => n2046);
   U2346 : NR2I port map( A => n2032, B => n4993, Z => n2128);
   U2348 : NR2I port map( A => v_RAM_OUT0_13_port, B => n1900, Z => n2367);
   U2349 : AO1P port map( A => n4998, B => n2306, C => n2369, D => n2370, Z => 
                           n2363);
   U2350 : NR2I port map( A => n2089_port, B => n4690, Z => n2370);
   U2351 : NR2I port map( A => n4955, B => n4970, Z => n2089_port);
   U2356 : ND2I port map( A => n4701, B => n2281, Z => n2227);
   U2359 : AO1P port map( A => n4360, B => n4982, C => n2378, D => n2379, Z => 
                           n2376);
   U2363 : ND2I port map( A => n1906, B => n2226, Z => n2261);
   U2364 : ND2I port map( A => n2186, B => n4391, Z => n2226);
   U2366 : AO1P port map( A => n4702, B => n4994, C => n2381, D => n2205, Z => 
                           n2375);
   U2368 : ND2I port map( A => n2281, B => n2153, Z => n2382);
   U2370 : ND2I port map( A => n2093, B => n2162, Z => n2067);
   U2371 : NR2I port map( A => n5069, B => n2095, Z => n2331);
   U2375 : ND2I port map( A => n2344, B => n2212, Z => n2038);
   U2377 : ND2I port map( A => n2178, B => n2162, Z => n2192);
   U2378 : NR2I port map( A => n4361, B => v_RAM_OUT0_13_port, Z => n2054);
   U2379 : NR2I port map( A => n4359, B => v_RAM_OUT0_13_port, Z => n2065);
   U2380 : NR2I port map( A => n4972, B => n4964, Z => n2386);
   U2382 : ND2I port map( A => n4977, B => v_RAM_OUT0_8_port, Z => n2162);
   U2383 : AO1P port map( A => n4360, B => n2064, C => n2387, D => n2241, Z => 
                           n2383);
   -- U2384 : ND2I port map( A => n2075, B => n4361, Z => n2241);--changing ND2I with NR2I
   U2384 : NR2I port map( A => n2075, B => n4361, Z => n2241);
   U2386 : ND2I port map( A => n4977, B => n2245, Z => n2166);
   U2387 : ND2I port map( A => v_RAM_OUT0_8_port, B => n2186, Z => n2245);
   U2391 : ND2I port map( A => n2390, B => n4529, Z => n2388);
   U2393 : ND2I port map( A => n2024, B => n4706, Z => n2020);
   U2394 : ND2I port map( A => n4706, B => n1602, Z => n2024);
   U2398 : AO1P port map( A => n4910, B => n2394, C => n1895, D => n2395, Z => 
                           n2393);
   U2404 : NR2I port map( A => n4976, B => n2095, Z => n1916);
   U2407 : NR2I port map( A => n4987, B => n4997, Z => n2402);
   U2410 : ND2I port map( A => n4378, B => n4516, Z => n1877);
   U2412 : ND2I port map( A => n2154, B => n2121, Z => n1907);
   U2413 : ND2I port map( A => v_RAM_OUT0_8_port, B => n2064, Z => n2154);
   U2415 : ND2I port map( A => n4360, B => n4516, Z => n2183);
   U2417 : ND2I port map( A => n4379, B => n4516, Z => n2318);
   U2419 : ND2I port map( A => v_RAM_OUT0_14_port, B => v_RAM_OUT0_8_port, Z =>
                           n1906);
   U2421 : ND2I port map( A => n1901, B => n2305, Z => n2404);
   U2422 : ND2I port map( A => n2121, B => n2167, Z => n2305);
   U2423 : ND2I port map( A => n4964, B => v_RAM_OUT0_8_port, Z => n2167);
   U2424 : ND2I port map( A => n4707, B => n4359, Z => n1901);
   U2425 : AO1P port map( A => n4989, B => v_RAM_OUT0_10_port, C => n2405, D =>
                           n2406, Z => n2403);
   U2427 : NR2I port map( A => n4983, B => n4997, Z => n2407);
   U2429 : ND2I port map( A => v_RAM_OUT0_8_port, B => n2408, Z => n2281);
   U2431 : ND2I port map( A => n4391, B => n2153, Z => n2075);
   U2433 : NR2I port map( A => n4960, B => n2061, Z => n2372);
   U2437 : ND2I port map( A => n2212, B => n2094, Z => n2190);
   U2438 : ND2I port map( A => v_RAM_OUT0_8_port, B => n4509, Z => n2094);
   U2439 : ND2I port map( A => n2306, B => n4391, Z => n2212);
   U2440 : ND2I port map( A => n1914, B => n2186, Z => n1913);
   U2441 : AO1P port map( A => n2410, B => n4906, C => n2411, D => n4908, Z => 
                           n1890);
   U2444 : ND2I port map( A => n2416, B => n2417, Z => n2415);
   U2447 : NR2I port map( A => n4960, B => n2095, Z => n2158);
   U2449 : ND2I port map( A => n4391, B => n4509, Z => n2072);
   U2451 : ND2I port map( A => n2344, B => n2121, Z => n2098);
   U2452 : ND2I port map( A => v_RAM_OUT0_14_port, B => n4391, Z => n2121);
   U2453 : ND2I port map( A => n4990, B => v_RAM_OUT0_8_port, Z => n2344);
   U2455 : ND2I port map( A => v_RAM_OUT0_14_port, B => n4412, Z => n2186);
   U2457 : ND2I port map( A => v_RAM_OUT0_13_port, B => v_RAM_OUT0_15_port, Z 
                           => n2074);
   U2461 : NR2I port map( A => n4970, B => n2061, Z => n2159);
   U2463 : ND2I port map( A => n4971, B => n4391, Z => n2178);
   U2467 : NR2I port map( A => n4976, B => n2061, Z => n1900);
   U2468 : NR2I port map( A => n4412, B => n4391, Z => n2061);
   U2470 : ND2I port map( A => n4977, B => n4391, Z => n2044);
   U2472 : ND2I port map( A => n4963, B => v_RAM_OUT0_10_port, Z => n2087_port)
                           ;
   U2474 : ND2I port map( A => n4964, B => n4391, Z => n2347);
   U2475 : ND2I port map( A => n2408, B => n1914, Z => n2144);
   U2477 : ND2I port map( A => v_RAM_OUT0_15_port, B => n4516, Z => n1912);
   U2478 : AO1P port map( A => n2093, B => n4379, C => n4691, D => n2419, Z => 
                           n2411);
   U2480 : ND2I port map( A => n2113, B => v_RAM_OUT0_10_port, Z => n1878);
   U2481 : NR2I port map( A => n2408, B => n4391, Z => n2113);
   U2482 : ND2I port map( A => n4701, B => n2215, Z => n2420);
   U2483 : NR2I port map( A => n4995, B => n2032, Z => n2215);
   U2484 : NR2I port map( A => n4391, B => v_RAM_OUT0_11_port, Z => n2032);
   U2486 : ND2I port map( A => n4391, B => n2408, Z => n2047);
   U2488 : NR2I port map( A => n2095, B => n4993, Z => n2380);
   U2490 : ND2I port map( A => n4994, B => n4391, Z => n2060);
   U2492 : NR2I port map( A => n2153, B => n4391, Z => n2095);
   U2493 : ND2I port map( A => v_RAM_OUT0_13_port, B => n4396, Z => n1898);
   U2494 : ND2I port map( A => n4391, B => n4412, Z => n2093);
   U2496 : ND2I port map( A => n4516, B => n4396, Z => n1897);
   U2500 : ND2I port map( A => n4964, B => n4379, Z => n2110);
   U2506 : NR2I port map( A => n4980, B => n4965, Z => n2234);
   U2508 : ND2I port map( A => n2064, B => n4391, Z => n2130);
   U2510 : ND2I port map( A => v_RAM_OUT0_11_port, B => n4509, Z => n2064);
   U2512 : ND2I port map( A => v_RAM_OUT0_8_port, B => n2153, Z => n1914);
   U2514 : ND2I port map( A => v_RAM_OUT0_10_port, B => n4404, Z => n2043);
   U2517 : ND2I port map( A => v_RAM_OUT0_8_port, B => n2306, Z => n2120);
   U2518 : ND2I port map( A => n2153, B => n2408, Z => n2306);
   U2519 : ND2I port map( A => v_RAM_OUT0_11_port, B => v_RAM_OUT0_14_port, Z 
                           => n2408);
   U2520 : ND2I port map( A => n4509, B => n4412, Z => n2153);
   U2527 : ND2I port map( A => n2425, B => n4435, Z => n2423);
   U2532 : ND2I port map( A => n2429, B => n4424, Z => n2427);
   -- U2538 : ND2I port map( A => n3840, B => n4655, Z => n423);--changing ND2I with EOI
   U2538 : EOI port map( A => n3840, B => n4655, Z => n423);
   U2542 : ND2I port map( A => n2433, B => n4557, Z => n2431);
   U2547 : ND2I port map( A => n2436, B => n4538, Z => n2434);
   U2551 : ND2I port map( A => n2440, B => n4537, Z => n2439);
   U2558 : ND2I port map( A => n2451, B => n2452, Z => n2450);
   U2563 : ND2I port map( A => n2462, B => n4556, Z => n2460);
   U2567 : ND2I port map( A => n2466, B => n4555, Z => n2465);
   U2571 : ND2I port map( A => n2426, B => n4706, Z => n2422);
   U2572 : ND2I port map( A => n4706, B => n1702, Z => n2426);
   U2586 : ND2I port map( A => n2494, B => n4593, Z => n2491);
   U2600 : NR2I port map( A => n4362, B => n4499, Z => n2525);
   U2609 : AO1P port map( A => n5043, B => n4914, C => n2547, D => n2548, Z => 
                           n2536);
   U2617 : ND2I port map( A => n2529, B => n2562, Z => n2509);
   U2624 : ND2I port map( A => n2572, B => n4428, Z => n2570);
   U2629 : AO1P port map( A => n2580, B => n4499, C => n2581, D => n2582, Z => 
                           n2579);
   U2632 : ND2I port map( A => n4875, B => n2589, Z => n2580);
   U2638 : ND2I port map( A => n4887, B => n4362, Z => n2600);
   U2641 : ND2I port map( A => n2605, B => n2606, Z => n2561);
   U2643 : ND2I port map( A => n2609, B => n2610, Z => n2574);
   U2645 : AO1P port map( A => n4357, B => n4912, C => n2615, D => n2616, Z => 
                           n2612);
   U2646 : NR2I port map( A => n1959, B => n2584, Z => n2616);
   U2649 : AO1P port map( A => n4703, B => n2621, C => n2622, D => n2623, Z => 
                           n2620);
   U2651 : NR2I port map( A => n4913, B => n4704, Z => n2622);
   U2657 : AO1P port map( A => n4372, B => n2632, C => n2633, D => n2634, Z => 
                           n2626);
   U2660 : ND2I port map( A => n2625, B => n1955, Z => n2632);
   U2664 : ND2I port map( A => n2638, B => n4413, Z => n2636);
   U2668 : NR2I port map( A => n2643, B => n2644, Z => n2642);
   U2678 : AO1P port map( A => n4703, B => n2559, C => v_RAM_OUT0_25_port, D =>
                           n2662, Z => n2661);
   U2679 : NR2I port map( A => n4704, B => n2617, Z => n2662);
   U2683 : NR2I port map( A => v_RAM_OUT0_28_port, B => n4871, Z => n2667);
   U2684 : ND2I port map( A => v_RAM_OUT0_31_port, B => n2670, Z => n2641);
   U2686 : AO1P port map( A => n4357, B => n2673, C => n2674, D => n2675, Z => 
                           n2672);
   U2689 : ND2I port map( A => n2583, B => n2542, Z => n2673);
   U2698 : AO1P port map( A => n4894, B => n4357, C => n2691, D => n2692, Z => 
                           n2679);
   U2700 : NR2I port map( A => n4883, B => n4894, Z => n2565);
   U2704 : ND2I port map( A => n2698, B => n4592, Z => n2695);
   U2706 : ND2I port map( A => n2699, B => n2700, Z => n1621);
   U2715 : ND2I port map( A => n2542, B => n2714, Z => n2684);
   U2716 : NR2I port map( A => n4892, B => n2715, Z => n2689);
   U2718 : NR2I port map( A => v_RAM_OUT0_29_port, B => n1959, Z => n2709);
   U2722 : ND2I port map( A => n2665, B => n2618, Z => n2706);
   U2726 : NR2I port map( A => n2721, B => n4704, Z => n2692);
   U2731 : NR2I port map( A => n4866, B => n4896, Z => n2729);
   U2738 : AO1P port map( A => n4357, B => n2735, C => n2736, D => n2737, Z => 
                           n2734);
   U2741 : ND2I port map( A => n2542, B => n2562, Z => n2735);
   U2748 : ND2I port map( A => n2745, B => n4443, Z => n2743);
   U2753 : ND2I port map( A => n2753, B => n2754, Z => n2752);
   U2758 : ND2I port map( A => n4372, B => n2665, Z => n2757);
   U2761 : ND2I port map( A => n4913, B => n2549, Z => n2568);
   U2765 : ND2I port map( A => n2529, B => n2739, Z => n2765);
   U2767 : ND2I port map( A => n2617, B => n2714, Z => n2768);
   U2768 : NR2I port map( A => n4912, B => n4898, Z => n2767);
   U2769 : NR2I port map( A => n4898, B => n4915, Z => n2762);
   U2772 : AO1P port map( A => n4703, B => n2688, C => n2773, D => n2774, Z => 
                           n2772);
   U2773 : NR2I port map( A => n4704, B => n2618, Z => n2774);
   U2775 : ND2I port map( A => n2507, B => n4895, Z => n2688);
   U2777 : AO1P port map( A => n4869, B => n4372, C => n2776, D => n2777, Z => 
                           n2771);
   U2780 : NR2I port map( A => n4887, B => n4893, Z => n2601);
   U2782 : AO1P port map( A => n4916, B => n5062, C => n2781, D => n2782, Z => 
                           n2779);
   U2783 : NR2I port map( A => n4898, B => n2783, Z => n2782);
   U2785 : AO1P port map( A => n1959, B => n2784, C => n1986, D => n4499, Z => 
                           n2781);
   U2786 : ND2I port map( A => n2785, B => n4362, Z => n2784);
   U2788 : ND2I port map( A => n2738, B => n2618, Z => n2785);
   U2789 : ND2I port map( A => n2617, B => n1955, Z => n2532);
   U2791 : ND2I port map( A => n2790, B => n4528, Z => n2789);
   U2801 : ND2I port map( A => n2529, B => n2676, Z => n2761);
   U2807 : ND2I port map( A => n2507, B => n2606, Z => n2802);
   U2809 : ND2I port map( A => n2803, B => n2605, Z => n2593);
   U2810 : NR2I port map( A => n4891, B => n4869, Z => n2755);
   U2813 : ND2I port map( A => n2586, B => n2713, Z => n2533);
   U2815 : NR2I port map( A => n2806, B => n2807, Z => n2793);
   U2818 : ND2I port map( A => n2759, B => n2583, Z => n2657);
   U2819 : NR2I port map( A => n4901, B => n4869, Z => n2742);
   U2823 : ND2I port map( A => n2811, B => n2812, Z => n2810);
   U2831 : ND2I port map( A => n4915, B => n4394, Z => n2606);
   U2833 : ND2I port map( A => n4703, B => n2584, Z => n2814);
   U2836 : ND2I port map( A => n4686, B => n2677, Z => n2821);
   U2837 : ND2I port map( A => v_RAM_OUT0_27_port, B => n4394, Z => n2677);
   U2839 : ND2I port map( A => n2625, B => n2618, Z => n2621);
   U2840 : AN2I port map( A => n2690, B => n2587, Z => n2707);
   U2846 : ND2I port map( A => n2826, B => n4442, Z => n2824);
   U2853 : ND2I port map( A => n2507, B => n2635, Z => n2608);
   U2857 : ND2I port map( A => n2690, B => n2586, Z => n2503);
   U2859 : ND2I port map( A => n2587, B => n2654, Z => n2719);
   U2860 : ND2I port map( A => n4703, B => n2708, Z => n2836);
   U2861 : ND2I port map( A => n2584, B => n2587, Z => n2708);
   U2864 : NR2I port map( A => n2590, B => n4891, Z => n1958);
   U2867 : ND2I port map( A => n2562, B => n2654, Z => n2523);
   U2869 : NR2I port map( A => n4913, B => n4898, Z => n2842);
   U2872 : NR2I port map( A => n2847, B => n2848, Z => n2846);
   U2874 : NR2I port map( A => n4882, B => n4899, Z => n2756);
   U2877 : AO1P port map( A => n4357, B => n2559, C => n2851, D => n2852, Z => 
                           n2845);
   U2880 : ND2I port map( A => n2676, B => n2665, Z => n2854);
   U2881 : NR2I port map( A => n4901, B => n4916, Z => n2853);
   U2883 : ND2I port map( A => n2529, B => n2587, Z => n2559);
   U2884 : ND2I port map( A => n4913, B => v_RAM_OUT0_24_port, Z => n2587);
   U2887 : ND2I port map( A => n2529, B => n4686, Z => n2860);
   U2888 : NR2I port map( A => n4914, B => n4891, Z => n2859);
   U2890 : ND2I port map( A => v_RAM_OUT0_24_port, B => n2550, Z => n2583);
   U2892 : ND2I port map( A => n2739, B => n2713, Z => n2850);
   U2893 : ND2I port map( A => n2550, B => n4394, Z => n2713);
   U2894 : NR2I port map( A => n1959, B => n4499, Z => n2527);
   U2895 : ND2I port map( A => n2714, B => n2635, Z => n2861);
   U2896 : ND2I port map( A => n4916, B => n4394, Z => n2635);
   U2898 : ND2I port map( A => n2690, B => n2605, Z => n2678);
   U2902 : ND2I port map( A => n2865, B => n4454, Z => n2864);
   U2906 : ND2I port map( A => n2495, B => n1527, Z => n2490);
   U2907 : ND2I port map( A => n1527, B => n1702, Z => n2495);
   U2913 : ND2I port map( A => n4499, B => n4410, Z => n1949);
   U2918 : ND2I port map( A => n4703, B => n2721, Z => n2872);
   U2919 : ND2I port map( A => n2624, B => n2654, Z => n2721);
   U2920 : ND2I port map( A => n4912, B => n4394, Z => n2654);
   U2924 : ND2I port map( A => n2562, B => n2690, Z => n2649);
   U2925 : ND2I port map( A => v_RAM_OUT0_24_port, B => n4508, Z => n2562);
   U2926 : ND2I port map( A => n4686, B => n2550, Z => n1988);
   U2927 : ND2I port map( A => n2617, B => n2605, Z => n1986);
   U2928 : ND2I port map( A => n4914, B => v_RAM_OUT0_24_port, Z => n2605);
   U2930 : ND2I port map( A => v_RAM_OUT0_25_port, B => n4410, Z => n1947);
   U2933 : ND2I port map( A => n2759, B => n4686, Z => n2619);
   U2936 : NR2I port map( A => n4881, B => n4893, Z => n2655);
   U2938 : ND2I port map( A => v_RAM_OUT0_24_port, B => v_RAM_OUT0_27_port, Z 
                           => n2624);
   U2940 : ND2I port map( A => n4394, B => n2665, Z => n2542);
   U2942 : NR2I port map( A => n2625, B => n4362, Z => n2874);
   U2943 : ND2I port map( A => n4914, B => n4394, Z => n2625);
   U2945 : ND2I port map( A => n2617, B => n2586, Z => n2552);
   U2946 : ND2I port map( A => n4915, B => v_RAM_OUT0_24_port, Z => n2586);
   U2948 : ND2I port map( A => v_RAM_OUT0_30_port, B => n4411, Z => n2550);
   U2949 : NR2I port map( A => n1959, B => v_RAM_OUT0_25_port, Z => n2522);
   U2950 : ND2I port map( A => n4898, B => n5063, Z => n2879);
   U2955 : NR2I port map( A => n4881, B => n4896, Z => n2591);
   U2957 : ND2I port map( A => n4508, B => n4394, Z => n2738);
   U2963 : ND2I port map( A => v_RAM_OUT0_29_port, B => n4499, Z => n2541);
   U2966 : NR2I port map( A => n4882, B => n4897, Z => n2652);
   U2969 : ND2I port map( A => n4394, B => n2759, Z => n2528);
   U2972 : ND2I port map( A => n4916, B => v_RAM_OUT0_24_port, Z => n1955);
   U2975 : ND2I port map( A => n4411, B => n4394, Z => n2529);
   U2978 : NR2I port map( A => n4896, B => n2715, Z => n1977);
   U2979 : NR2I port map( A => n2590, B => v_RAM_OUT0_24_port, Z => n2715);
   U2981 : ND2I port map( A => n4912, B => v_RAM_OUT0_24_port, Z => n2714);
   U2983 : ND2I port map( A => n2507, B => n2690, Z => n2540);
   U2984 : ND2I port map( A => n2590, B => n4394, Z => n2690);
   U2985 : ND2I port map( A => v_RAM_OUT0_24_port, B => n4411, Z => n2507);
   U2987 : ND2I port map( A => n4704, B => n1959, Z => n1978);
   U2989 : ND2I port map( A => v_RAM_OUT0_25_port, B => v_RAM_OUT0_29_port, Z 
                           => n2544);
   U2992 : ND2I port map( A => v_RAM_OUT0_24_port, B => n2590, Z => n2618);
   U2993 : ND2I port map( A => n2665, B => n2759, Z => n2590);
   U2994 : NR2I port map( A => n4687, B => v_RAM_OUT0_25_port, Z => n2531);
   U2996 : ND2I port map( A => n4372, B => n4499, Z => n2519);
   U2999 : ND2I port map( A => n2676, B => n2617, Z => n2808);
   U3000 : ND2I port map( A => v_RAM_OUT0_24_port, B => n2759, Z => n2676);
   U3001 : ND2I port map( A => v_RAM_OUT0_27_port, B => v_RAM_OUT0_30_port, Z 
                           => n2759);
   U3003 : ND2I port map( A => n4357, B => v_RAM_OUT0_25_port, Z => n2534);
   U3007 : ND2I port map( A => n4372, B => v_RAM_OUT0_25_port, Z => n2530);
   U3011 : ND2I port map( A => v_RAM_OUT0_24_port, B => v_RAM_OUT0_30_port, Z 
                           => n2739);
   U3012 : ND2I port map( A => n4703, B => n2728, Z => n2890);
   U3013 : ND2I port map( A => n4686, B => n2803, Z => n2728);
   U3014 : ND2I port map( A => n2584, B => n4394, Z => n2803);
   U3015 : ND2I port map( A => v_RAM_OUT0_24_port, B => n2665, Z => n1973);
   U3016 : ND2I port map( A => n4508, B => n4411, Z => n2665);
   U3018 : ND2I port map( A => n4362, B => n4368, Z => n1959);
   U3021 : ND2I port map( A => n2549, B => n2617, Z => n2822);
   U3024 : ND2I port map( A => v_RAM_OUT0_24_port, B => n2584, Z => n2549);
   U3028 : ND2I port map( A => n4371, B => v_RAM_OUT0_25_port, Z => n2585);
   U3031 : ND2I port map( A => n4371, B => n4499, Z => n2651);
   U3039 : ND2I port map( A => n2896, B => n4522, Z => n2894);
   U3054 : NR2I port map( A => n4365, B => n4498, Z => n2930);
   U3062 : AO1P port map( A => n5038, B => n4925, C => n2951, D => n2952, Z => 
                           n2942);
   U3070 : ND2I port map( A => n2935, B => n2965, Z => n2913);
   U3077 : ND2I port map( A => n2974, B => n4609, Z => n2971);
   U3083 : AO1P port map( A => n2983, B => n4498, C => n2984, D => n2985, Z => 
                           n2982);
   U3086 : ND2I port map( A => n4931, B => n2992, Z => n2983);
   U3092 : ND2I port map( A => n4928, B => n4365, Z => n3002);
   U3095 : ND2I port map( A => n3008, B => n3009, Z => n2964);
   U3097 : ND2I port map( A => n3012, B => n3013, Z => n2976);
   U3099 : AO1P port map( A => n4355, B => n4935, C => n3017, D => n3018, Z => 
                           n3014);
   U3100 : NR2I port map( A => n2957, B => n2987, Z => n3018);
   U3103 : AO1P port map( A => n4699, B => n3024, C => n3025, D => n3026, Z => 
                           n3023);
   U3105 : NR2I port map( A => n4937, B => n4698, Z => n3025);
   U3111 : AO1P port map( A => n4374, B => n3036, C => n3037, D => n3038, Z => 
                           n3030);
   U3114 : ND2I port map( A => n3028, B => n3007, Z => n3036);
   U3118 : ND2I port map( A => n3042, B => n4521, Z => n3040);
   U3123 : NR2I port map( A => n3047, B => n3048, Z => n3046);
   U3133 : AO1P port map( A => n4699, B => n2962, C => v_RAM_OUT0_17_port, D =>
                           n3067, Z => n3066);
   U3134 : NR2I port map( A => n4698, B => n3019, Z => n3067);
   U3138 : NR2I port map( A => v_RAM_OUT0_20_port, B => n4947, Z => n3072);
   U3139 : ND2I port map( A => v_RAM_OUT0_23_port, B => n3075, Z => n3045);
   U3141 : AO1P port map( A => n4355, B => n3078, C => n3079, D => n3080, Z => 
                           n3077);
   U3144 : ND2I port map( A => n2986, B => n2947, Z => n3078);
   U3153 : AO1P port map( A => n4951, B => n4355, C => n3096, D => n3097, Z => 
                           n3084);
   U3155 : NR2I port map( A => n5065, B => n4951, Z => n2968);
   U3159 : ND2I port map( A => n3103, B => n4608, Z => n3100);
   U3162 : ND2I port map( A => n3104, B => n3105, Z => n1661);
   U3171 : ND2I port map( A => n2947, B => n3118, Z => n3089);
   U3172 : NR2I port map( A => n4917, B => n3119, Z => n3094);
   U3174 : NR2I port map( A => v_RAM_OUT0_21_port, B => n2957, Z => n3114);
   U3178 : ND2I port map( A => n3070, B => n3020, Z => n3111);
   U3182 : NR2I port map( A => n3125, B => n4698, Z => n3097);
   U3188 : NR2I port map( A => n4945, B => n4934, Z => n3133);
   U3195 : AO1P port map( A => n4355, B => n3139, C => n3140, D => n3141, Z => 
                           n3138);
   U3198 : ND2I port map( A => n2947, B => n2965, Z => n3139);
   U3205 : ND2I port map( A => n3149, B => n4536, Z => n3147);
   U3211 : ND2I port map( A => n3157, B => n3158, Z => n3156);
   U3216 : ND2I port map( A => n4374, B => n3070, Z => n3161);
   U3219 : ND2I port map( A => n4937, B => n2953, Z => n2970);
   U3223 : ND2I port map( A => n2935, B => n3143, Z => n3169);
   U3225 : ND2I port map( A => n3019, B => n3118, Z => n3172);
   U3226 : NR2I port map( A => n4935, B => n4953, Z => n3171);
   U3227 : NR2I port map( A => n4953, B => n4946, Z => n3166);
   U3230 : AO1P port map( A => n4699, B => n3093, C => n3177, D => n3178, Z => 
                           n3176);
   U3231 : NR2I port map( A => n4698, B => n3020, Z => n3178);
   U3233 : ND2I port map( A => n2911, B => n4939, Z => n3093);
   U3235 : AO1P port map( A => n5067, B => n4374, C => n3180, D => n3181, Z => 
                           n3175);
   U3238 : NR2I port map( A => n4928, B => n5068, Z => n3003);
   U3240 : AO1P port map( A => n4952, B => n5054, C => n3186, D => n3187, Z => 
                           n3184);
   U3241 : NR2I port map( A => n4953, B => n3188, Z => n3187);
   U3243 : AO1P port map( A => n2957, B => n3189, C => n1710, D => n4498, Z => 
                           n3186);
   U3244 : ND2I port map( A => n3190, B => n4365, Z => n3189);
   U3246 : ND2I port map( A => n3142, B => n3020, Z => n3190);
   U3250 : ND2I port map( A => n3194, B => n4535, Z => n3192);
   U3256 : AO1P port map( A => n4937, B => n1687, C => n3198, D => n3199, Z => 
                           n3197);
   U3257 : NR2I port map( A => n4700, B => n3007, Z => n3199);
   U3260 : ND2I port map( A => n3019, B => n3007, Z => n3182);
   U3267 : ND2I port map( A => n4699, B => n2987, Z => n3201);
   U3270 : ND2I port map( A => n4683, B => n3082, Z => n3207);
   U3272 : ND2I port map( A => n3028, B => n3020, Z => n3024);
   U3273 : AN2I port map( A => n3095, B => n2990, Z => n3112);
   U3281 : ND2I port map( A => n2935, B => n3081, Z => n3165);
   U3287 : ND2I port map( A => n2911, B => n3009, Z => n3220);
   U3288 : ND2I port map( A => n4946, B => n4393, Z => n3009);
   U3290 : ND2I port map( A => n3221, B => n3008, Z => n2995);
   U3291 : NR2I port map( A => n4948, B => n5067, Z => n3159);
   U3293 : ND2I port map( A => v_RAM_OUT0_21_port, B => n4498, Z => n2946);
   U3296 : ND2I port map( A => n2989, B => n3117, Z => n2939);
   U3298 : ND2I port map( A => v_RAM_OUT0_17_port, B => v_RAM_OUT0_21_port, Z 
                           => n2949);
   U3299 : NR2I port map( A => n3225, B => n3226, Z => n3211);
   U3302 : ND2I port map( A => n3163, B => n2986, Z => n3062);
   U3303 : NR2I port map( A => n4926, B => n5067, Z => n3146);
   U3305 : ND2I port map( A => v_RAM_OUT0_19_port, B => n4393, Z => n3082);
   U3309 : ND2I port map( A => n3230, B => n4567, Z => n3228);
   U3317 : ND2I port map( A => n2911, B => n3039, Z => n3011);
   U3322 : ND2I port map( A => n3095, B => n2989, Z => n2907);
   U3324 : ND2I port map( A => n2990, B => n3058, Z => n3123);
   U3325 : ND2I port map( A => n4699, B => n3113, Z => n3240);
   U3326 : ND2I port map( A => n2987, B => n2990, Z => n3113);
   U3330 : NR2I port map( A => n1688, B => n4948, Z => n1689);
   U3333 : ND2I port map( A => n2965, B => n3058, Z => n2927);
   U3335 : NR2I port map( A => n4937, B => n4953, Z => n3246);
   U3338 : NR2I port map( A => n3251, B => n3252, Z => n3250);
   U3340 : NR2I port map( A => n4954, B => n4943, Z => n3160);
   U3343 : AO1P port map( A => n4355, B => n2962, C => n3255, D => n3256, Z => 
                           n3249);
   U3346 : ND2I port map( A => n3081, B => n3070, Z => n3258);
   U3347 : NR2I port map( A => n4926, B => n4952, Z => n3257);
   U3349 : ND2I port map( A => n2935, B => n2990, Z => n2962);
   U3350 : ND2I port map( A => n4937, B => v_RAM_OUT0_16_port, Z => n2990);
   U3353 : ND2I port map( A => n2935, B => n4683, Z => n3264);
   U3354 : NR2I port map( A => n4925, B => n4948, Z => n3263);
   U3356 : ND2I port map( A => v_RAM_OUT0_16_port, B => n2954, Z => n2986);
   U3358 : ND2I port map( A => n3143, B => n3117, Z => n3254);
   U3359 : ND2I port map( A => n2954, B => n4393, Z => n3117);
   U3360 : NR2I port map( A => n2957, B => n4498, Z => n2932);
   U3361 : ND2I port map( A => n3118, B => n3039, Z => n3265);
   U3362 : ND2I port map( A => n4952, B => n4393, Z => n3039);
   U3364 : ND2I port map( A => n3095, B => n3008, Z => n3083);
   U3370 : ND2I port map( A => n3268, B => n4534, Z => n3266);
   U3373 : ND2I port map( A => n2897, B => n1527, Z => n2893);
   U3374 : ND2I port map( A => n1527, B => n1754, Z => n2897);
   U3381 : ND2I port map( A => n3081, B => n3019, Z => n3227);
   U3383 : ND2I port map( A => v_RAM_OUT0_16_port, B => v_RAM_OUT0_22_port, Z 
                           => n3143);
   U3384 : ND2I port map( A => n4699, B => n3132, Z => n3274);
   U3385 : ND2I port map( A => n4683, B => n3221, Z => n3132);
   U3386 : ND2I port map( A => n2987, B => n4393, Z => n3221);
   U3388 : ND2I port map( A => n2953, B => n3019, Z => n3208);
   U3389 : ND2I port map( A => v_RAM_OUT0_16_port, B => n2987, Z => n2953);
   U3390 : AO1P port map( A => n5056, B => n4683, C => n3277, D => n3278, Z => 
                           n3272);
   U3391 : AN2I port map( A => n5053, B => n1725, Z => n3278);
   U3392 : NR2I port map( A => n4934, B => n3119, Z => n1725);
   U3393 : NR2I port map( A => n1688, B => v_RAM_OUT0_16_port, Z => n3119);
   U3396 : ND2I port map( A => n4369, B => v_RAM_OUT0_17_port, Z => n2988);
   U3400 : NR2I port map( A => n4954, B => n5066, Z => n3056);
   U3403 : ND2I port map( A => n4393, B => n3163, Z => n2933);
   U3406 : ND2I port map( A => n4952, B => v_RAM_OUT0_16_port, Z => n3007);
   U3409 : ND2I port map( A => n4406, B => n4393, Z => n2935);
   U3413 : ND2I port map( A => v_RAM_OUT0_17_port, B => n4409, Z => n2906);
   U3417 : ND2I port map( A => n2965, B => n3095, Z => n3053);
   U3418 : ND2I port map( A => v_RAM_OUT0_16_port, B => n4501, Z => n2965);
   U3419 : ND2I port map( A => n4683, B => n2954, Z => n1713);
   U3420 : ND2I port map( A => n3019, B => n3008, Z => n1710);
   U3421 : ND2I port map( A => n4925, B => v_RAM_OUT0_16_port, Z => n3008);
   U3422 : ND2I port map( A => n4698, B => n2957, Z => n1712);
   U3423 : ND2I port map( A => n4498, B => n4409, Z => n2904);
   U3429 : ND2I port map( A => n2911, B => n3095, Z => n1722);
   U3430 : ND2I port map( A => n1688, B => n4393, Z => n3095);
   U3431 : ND2I port map( A => v_RAM_OUT0_16_port, B => n4406, Z => n2911);
   U3432 : ND2I port map( A => n4699, B => n3125, Z => n3286);
   U3433 : ND2I port map( A => n3027, B => n3058, Z => n3125);
   U3434 : ND2I port map( A => n4935, B => n4393, Z => n3058);
   U3438 : ND2I port map( A => n4374, B => n4498, Z => n2923);
   U3439 : ND2I port map( A => n3163, B => n4683, Z => n3022);
   U3440 : ND2I port map( A => v_RAM_OUT0_16_port, B => n3070, Z => n1724);
   U3443 : NR2I port map( A => n4942, B => n5068, Z => n3060);
   U3445 : ND2I port map( A => v_RAM_OUT0_16_port, B => v_RAM_OUT0_19_port, Z 
                           => n3027);
   U3447 : ND2I port map( A => n4393, B => n3070, Z => n2947);
   U3449 : NR2I port map( A => n3028, B => n4365, Z => n3288);
   U3450 : ND2I port map( A => n4925, B => n4393, Z => n3028);
   U3454 : ND2I port map( A => n3019, B => n2989, Z => n2955);
   U3455 : ND2I port map( A => n4946, B => v_RAM_OUT0_16_port, Z => n2989);
   U3457 : ND2I port map( A => v_RAM_OUT0_22_port, B => n4406, Z => n2954);
   U3459 : NR2I port map( A => n2957, B => v_RAM_OUT0_17_port, Z => n2926);
   U3460 : ND2I port map( A => n4365, B => n4364, Z => n2957);
   U3461 : ND2I port map( A => v_RAM_OUT0_16_port, B => n1688, Z => n3020);
   U3463 : ND2I port map( A => n4355, B => v_RAM_OUT0_17_port, Z => n2940);
   U3465 : ND2I port map( A => n4953, B => n5055, Z => n3290);
   U3467 : ND2I port map( A => n4374, B => v_RAM_OUT0_17_port, Z => n2936);
   U3471 : ND2I port map( A => v_RAM_OUT0_16_port, B => n3163, Z => n3081);
   U3474 : ND2I port map( A => n3070, B => n3163, Z => n1688);
   U3475 : ND2I port map( A => v_RAM_OUT0_19_port, B => v_RAM_OUT0_22_port, Z 
                           => n3163);
   U3477 : ND2I port map( A => n4369, B => n4498, Z => n3055);
   U3483 : NR2I port map( A => n4942, B => n4934, Z => n2993);
   U3485 : ND2I port map( A => n4935, B => v_RAM_OUT0_16_port, Z => n3118);
   U3487 : ND2I port map( A => n4501, B => n4406, Z => n3070);
   U3490 : ND2I port map( A => n4501, B => n4393, Z => n3142);
   U3493 : NR2I port map( A => n4682, B => v_RAM_OUT0_17_port, Z => n2938);
   U3499 : ND2I port map( A => n3298, B => n4417, Z => n3296);
   U3513 : NR2I port map( A => n4363, B => n4497, Z => n3332);
   U3521 : AO1P port map( A => n5045, B => n5007, C => n3353, D => n3354, Z => 
                           n3344);
   U3529 : ND2I port map( A => n3337, B => n3367, Z => n3315);
   U3536 : ND2I port map( A => n3375, B => n4416, Z => n3373);
   U3541 : AO1P port map( A => n3384, B => n4497, C => n3385, D => n3386, Z => 
                           n3383);
   U3544 : ND2I port map( A => n5013, B => n3393, Z => n3384);
   U3550 : ND2I port map( A => n5010, B => n4363, Z => n3403);
   U3553 : ND2I port map( A => n3409, B => n3410, Z => n3366);
   U3555 : ND2I port map( A => n3413, B => n3414, Z => n3377);
   U3557 : AO1P port map( A => n4356, B => n5017, C => n3418, D => n3419, Z => 
                           n3415);
   U3558 : NR2I port map( A => n3359, B => n3388, Z => n3419);
   U3561 : AO1P port map( A => n4696, B => n3425, C => n3426, D => n3427, Z => 
                           n3424);
   U3563 : NR2I port map( A => n5019, B => n4695, Z => n3426);
   U3569 : AO1P port map( A => n4373, B => n3437, C => n3438, D => n3439, Z => 
                           n3431);
   U3572 : ND2I port map( A => n3429, B => n3408, Z => n3437);
   U3576 : ND2I port map( A => n3444, B => n4604, Z => n3441);
   U3580 : NR2I port map( A => n3449, B => n3450, Z => n3448);
   U3590 : AO1P port map( A => n4696, B => n3364, C => v_RAM_OUT0_1_port, D => 
                           n3469, Z => n3468);
   U3591 : NR2I port map( A => n4695, B => n3420, Z => n3469);
   U3595 : NR2I port map( A => v_RAM_OUT0_4_port, B => n5029, Z => n3474);
   U3596 : ND2I port map( A => v_RAM_OUT0_7_port, B => n3477, Z => n3447);
   U3598 : AO1P port map( A => n4356, B => n3480, C => n3481, D => n3482, Z => 
                           n3479);
   U3601 : ND2I port map( A => n3387, B => n3349, Z => n3480);
   U3610 : AO1P port map( A => n5033, B => n4356, C => n3498, D => n3499, Z => 
                           n3486);
   U3612 : NR2I port map( A => n5070, B => n5033, Z => n3370);
   U3616 : ND2I port map( A => n3504, B => n4547, Z => n3502);
   U3618 : ND2I port map( A => n3505, B => n3506, Z => n1581);
   U3627 : ND2I port map( A => n3349, B => n3519, Z => n3491);
   U3628 : NR2I port map( A => n4999, B => n3520, Z => n3496);
   U3630 : NR2I port map( A => v_RAM_OUT0_5_port, B => n3359, Z => n3515);
   U3634 : ND2I port map( A => n3472, B => n3421, Z => n3512);
   U3638 : NR2I port map( A => n3526, B => n4695, Z => n3499);
   U3644 : NR2I port map( A => n5027, B => n5016, Z => n3534);
   U3651 : AO1P port map( A => n4356, B => n3540, C => n3541, D => n3542, Z => 
                           n3539);
   U3654 : ND2I port map( A => n3349, B => n3367, Z => n3540);
   U3661 : ND2I port map( A => n3550, B => n4546, Z => n3548);
   U3666 : ND2I port map( A => n3558, B => n3559, Z => n3557);
   U3671 : ND2I port map( A => n4373, B => n3472, Z => n3562);
   U3674 : ND2I port map( A => n5019, B => n3355, Z => n3372);
   U3678 : ND2I port map( A => n3337, B => n3544, Z => n3570);
   U3680 : ND2I port map( A => n3420, B => n3519, Z => n3573);
   U3681 : NR2I port map( A => n5017, B => n5035, Z => n3572);
   U3682 : NR2I port map( A => n5035, B => n5028, Z => n3567);
   U3685 : AO1P port map( A => n4696, B => n3495, C => n3578, D => n3579, Z => 
                           n3577);
   U3686 : NR2I port map( A => n4695, B => n3421, Z => n3579);
   U3688 : ND2I port map( A => n3313, B => n5021, Z => n3495);
   U3690 : AO1P port map( A => n5072, B => n4373, C => n3581, D => n3582, Z => 
                           n3576);
   U3693 : NR2I port map( A => n5010, B => n5073, Z => n3404);
   U3695 : AO1P port map( A => n5034, B => n5048, C => n3587, D => n3588, Z => 
                           n3585);
   U3696 : NR2I port map( A => n5035, B => n3589, Z => n3588);
   U3698 : AO1P port map( A => n3359, B => n3590, C => n2474, D => n4497, Z => 
                           n3587);
   U3699 : ND2I port map( A => n3591, B => n4363, Z => n3590);
   U3701 : ND2I port map( A => n3543, B => n3421, Z => n3591);
   U3705 : ND2I port map( A => n3595, B => n4517, Z => n3593);
   U3710 : AO1P port map( A => n5019, B => n2453, C => n3599, D => n3600, Z => 
                           n3598);
   U3711 : NR2I port map( A => n4697, B => n3408, Z => n3600);
   U3714 : ND2I port map( A => n3420, B => n3408, Z => n3583);
   U3721 : ND2I port map( A => n4696, B => n3388, Z => n3602);
   U3724 : ND2I port map( A => n4679, B => n3484, Z => n3608);
   U3726 : ND2I port map( A => n3429, B => n3421, Z => n3425);
   U3727 : AN2I port map( A => n3497, B => n3391, Z => n3513);
   U3735 : ND2I port map( A => n3337, B => n3483, Z => n3566);
   U3741 : ND2I port map( A => n3313, B => n3410, Z => n3621);
   U3742 : ND2I port map( A => n5028, B => n4392, Z => n3410);
   U3744 : ND2I port map( A => n3622, B => n3409, Z => n3396);
   U3745 : NR2I port map( A => n5030, B => n5072, Z => n3560);
   U3747 : ND2I port map( A => v_RAM_OUT0_5_port, B => n4497, Z => n3348);
   U3750 : ND2I port map( A => n3390, B => n3518, Z => n3341);
   U3752 : ND2I port map( A => v_RAM_OUT0_1_port, B => v_RAM_OUT0_5_port, Z => 
                           n3351);
   U3753 : NR2I port map( A => n3626, B => n3627, Z => n3612);
   U3756 : ND2I port map( A => n3564, B => n3387, Z => n3464);
   U3757 : NR2I port map( A => n5008, B => n5072, Z => n3547);
   U3759 : ND2I port map( A => v_RAM_OUT0_3_port, B => n4392, Z => n3484);
   U3763 : ND2I port map( A => n3632, B => n4603, Z => n3629);
   U3770 : ND2I port map( A => n3313, B => n3440, Z => n3412);
   U3775 : ND2I port map( A => n3497, B => n3390, Z => n3309);
   U3777 : ND2I port map( A => n3391, B => n3460, Z => n3524);
   U3778 : ND2I port map( A => n4696, B => n3514, Z => n3642);
   U3779 : ND2I port map( A => n3388, B => n3391, Z => n3514);
   U3783 : NR2I port map( A => n2454, B => n5030, Z => n2455);
   U3786 : ND2I port map( A => n3367, B => n3460, Z => n3329);
   U3788 : NR2I port map( A => n5019, B => n5035, Z => n3648);
   U3791 : NR2I port map( A => n3653, B => n3654, Z => n3652);
   U3793 : NR2I port map( A => n5036, B => n5025, Z => n3561);
   U3796 : AO1P port map( A => n4356, B => n3364, C => n3657, D => n3658, Z => 
                           n3651);
   U3799 : ND2I port map( A => n3483, B => n3472, Z => n3660);
   U3800 : NR2I port map( A => n5008, B => n5034, Z => n3659);
   U3802 : ND2I port map( A => n3337, B => n3391, Z => n3364);
   U3803 : ND2I port map( A => n5019, B => v_RAM_OUT0_0_port, Z => n3391);
   U3806 : ND2I port map( A => n3337, B => n4679, Z => n3666);
   U3807 : NR2I port map( A => n5007, B => n5030, Z => n3665);
   U3809 : ND2I port map( A => v_RAM_OUT0_0_port, B => n3356, Z => n3387);
   U3811 : ND2I port map( A => n3544, B => n3518, Z => n3656);
   U3812 : ND2I port map( A => n3356, B => n4392, Z => n3518);
   U3813 : NR2I port map( A => n3359, B => n4497, Z => n3334);
   U3814 : ND2I port map( A => n3519, B => n3440, Z => n3667);
   U3815 : ND2I port map( A => n5034, B => n4392, Z => n3440);
   U3817 : ND2I port map( A => n3497, B => n3409, Z => n3485);
   U3823 : ND2I port map( A => n3670, B => n4545, Z => n3668);
   U3825 : ND2I port map( A => n3299, B => n4352, Z => n3295);
   U3826 : ND2I port map( A => n4352, B => n1754, Z => n3299);
   U3827 : ND2I port map( A => n3671, B => n4579, Z => n1754);
   U3836 : ND2I port map( A => n3483, B => n3420, Z => n3628);
   U3838 : ND2I port map( A => v_RAM_OUT0_0_port, B => v_RAM_OUT0_6_port, Z => 
                           n3544);
   U3839 : ND2I port map( A => n4696, B => n3533, Z => n3678);
   U3840 : ND2I port map( A => n4679, B => n3622, Z => n3533);
   U3841 : ND2I port map( A => n3388, B => n4392, Z => n3622);
   U3843 : ND2I port map( A => n3355, B => n3420, Z => n3609);
   U3844 : ND2I port map( A => v_RAM_OUT0_0_port, B => n3388, Z => n3355);
   U3845 : AO1P port map( A => n5050, B => n4679, C => n3681, D => n3682, Z => 
                           n3676);
   U3846 : AN2I port map( A => n5047, B => n2489, Z => n3682);
   U3847 : NR2I port map( A => n5016, B => n3520, Z => n2489);
   U3848 : NR2I port map( A => n2454, B => v_RAM_OUT0_0_port, Z => n3520);
   U3851 : ND2I port map( A => n4370, B => v_RAM_OUT0_1_port, Z => n3389);
   U3855 : NR2I port map( A => n5036, B => n5071, Z => n3458);
   U3858 : ND2I port map( A => n4392, B => n3564, Z => n3335);
   U3861 : ND2I port map( A => n5034, B => v_RAM_OUT0_0_port, Z => n3408);
   U3864 : ND2I port map( A => n4405, B => n4392, Z => n3337);
   U3868 : ND2I port map( A => v_RAM_OUT0_1_port, B => n4408, Z => n3308);
   U3872 : ND2I port map( A => n3367, B => n3497, Z => n3455);
   U3873 : ND2I port map( A => v_RAM_OUT0_0_port, B => n4500, Z => n3367);
   U3874 : ND2I port map( A => n4679, B => n3356, Z => n2477);
   U3875 : ND2I port map( A => n3420, B => n3409, Z => n2474);
   U3876 : ND2I port map( A => n5007, B => v_RAM_OUT0_0_port, Z => n3409);
   U3877 : ND2I port map( A => n4695, B => n3359, Z => n2476);
   U3878 : ND2I port map( A => n4497, B => n4408, Z => n3306);
   U3884 : ND2I port map( A => n3313, B => n3497, Z => n2486);
   U3885 : ND2I port map( A => n2454, B => n4392, Z => n3497);
   U3886 : ND2I port map( A => v_RAM_OUT0_0_port, B => n4405, Z => n3313);
   U3887 : ND2I port map( A => n4696, B => n3526, Z => n3690);
   U3888 : ND2I port map( A => n3428, B => n3460, Z => n3526);
   U3889 : ND2I port map( A => n5017, B => n4392, Z => n3460);
   U3893 : ND2I port map( A => n4373, B => n4497, Z => n3325);
   U3894 : ND2I port map( A => n3564, B => n4679, Z => n3423);
   U3895 : ND2I port map( A => v_RAM_OUT0_0_port, B => n3472, Z => n2488);
   U3898 : NR2I port map( A => n5024, B => n5073, Z => n3462);
   U3900 : ND2I port map( A => v_RAM_OUT0_0_port, B => v_RAM_OUT0_3_port, Z => 
                           n3428);
   U3902 : ND2I port map( A => n4392, B => n3472, Z => n3349);
   U3904 : NR2I port map( A => n3429, B => n4363, Z => n3692);
   U3905 : ND2I port map( A => n5007, B => n4392, Z => n3429);
   U3909 : ND2I port map( A => n3420, B => n3390, Z => n3357);
   U3910 : ND2I port map( A => n5028, B => v_RAM_OUT0_0_port, Z => n3390);
   U3912 : ND2I port map( A => v_RAM_OUT0_6_port, B => n4405, Z => n3356);
   U3914 : NR2I port map( A => n3359, B => v_RAM_OUT0_1_port, Z => n3328);
   U3915 : ND2I port map( A => n4363, B => n4367, Z => n3359);
   U3916 : ND2I port map( A => v_RAM_OUT0_0_port, B => n2454, Z => n3421);
   U3918 : ND2I port map( A => n4356, B => v_RAM_OUT0_1_port, Z => n3342);
   U3920 : ND2I port map( A => n5035, B => n5049, Z => n3694);
   U3922 : ND2I port map( A => n4373, B => v_RAM_OUT0_1_port, Z => n3338);
   U3926 : ND2I port map( A => v_RAM_OUT0_0_port, B => n3564, Z => n3483);
   U3929 : ND2I port map( A => n3472, B => n3564, Z => n2454);
   U3930 : ND2I port map( A => v_RAM_OUT0_3_port, B => v_RAM_OUT0_6_port, Z => 
                           n3564);
   U3932 : ND2I port map( A => n4370, B => n4497, Z => n3457);
   U3938 : NR2I port map( A => n5024, B => n5016, Z => n3394);
   U3940 : ND2I port map( A => n5017, B => v_RAM_OUT0_0_port, Z => n3519);
   U3942 : ND2I port map( A => n4500, B => n4405, Z => n3472);
   U3945 : ND2I port map( A => n4500, B => n4392, Z => n3543);
   U3948 : NR2I port map( A => n4678, B => v_RAM_OUT0_1_port, Z => n3340);
   U3952 : ND2I port map( A => n4677, B => n3699, Z => N192);
   U3955 : ND2I port map( A => n1425, B => n4395, Z => n1427);
   U3957 : NR2I port map( A => n4426, B => n4840, Z => n1425);
   U3959 : ND2I port map( A => n3700, B => n3701, Z => n4311);
   U3963 : ND2I port map( A => n3951, B => n1474, Z => n1481);
   U3967 : NR2I port map( A => n4713, B => RESET_I, Z => n3704);
   U3975 : AO1P port map( A => n1517, B => n4591, C => n3716, D => n3717, Z => 
                           n3715);
   U3997 : AO1P port map( A => n1517, B => n4427, C => n3728, D => n3729, Z => 
                           n3727);
   U4019 : AO1P port map( A => n1517, B => n4507, C => n3739, D => n3740, Z => 
                           n3738);
   U4041 : AO1P port map( A => n1517, B => n4590, C => n3750, D => n3751, Z => 
                           n3749);
   U4063 : AO1P port map( A => n1517, B => n4453, C => n3761, D => n3762, Z => 
                           n3760);
   U4085 : AO1P port map( A => n1517, B => n4544, C => n3772, D => n3773, Z => 
                           n3771);
   U4107 : AO1P port map( A => n1517, B => n4543, C => n3783, D => n3784, Z => 
                           n3782);
   U4127 : ND2I port map( A => n4366, B => n1354, Z => n1527);
   U4128 : AN2I port map( A => n1391, B => n4601, Z => n1354);
   U4132 : ND2I port map( A => n4366, B => n1351, Z => n1609);
   U4135 : AO1P port map( A => n1517, B => n4440, C => n3794, D => n3795, Z => 
                           n3793);
   U4137 : ND2I port map( A => n3796, B => n4862, Z => n1520);
   U4138 : ND2I port map( A => n2019, B => n4862, Z => n1521);
   U4143 : NR2I port map( A => n2391, B => n3800, Z => n1515);
   U4145 : NR2I port map( A => n3800, B => n2866, Z => n1516);
   U4147 : NR2I port map( A => n3798, B => n2391, Z => n1517);
   U4150 : ND2I port map( A => n3802, B => n2019, Z => n1510);
   U4151 : ND2I port map( A => n2019, B => n3803, Z => n1511);
   U4152 : NR2I port map( A => n4601, B => v_CALCULATION_CNTR_2_port, Z => 
                           n2019);
   U4154 : NR2I port map( A => n4861, B => n2866, Z => n1513);
   U4157 : AN2I port map( A => n3796, B => n3803, Z => n1508);
   U4159 : NR2I port map( A => n3798, B => n2866, Z => n1506);
   U4160 : ND2I port map( A => v_CALCULATION_CNTR_0_port, B => 
                           v_CALCULATION_CNTR_2_port, Z => n2866);
   U4161 : ND2I port map( A => v_CALCULATION_CNTR_3_port, B => n4863, Z => 
                           n3798);
   U4166 : ND2I port map( A => n3802, B => n3796, Z => n1509);
   U4167 : NR2I port map( A => v_CALCULATION_CNTR_2_port, B => 
                           v_CALCULATION_CNTR_0_port, Z => n3796);
   U4169 : NR2I port map( A => n4861, B => n2391, Z => n1507);
   U4173 : ND2I port map( A => n4407, B => n4384, Z => n2392);
   U4176 : ND2I port map( A => n1391, B => v_CALCULATION_CNTR_0_port, Z => 
                           n1485);
   U4177 : NR2I port map( A => n3800, B => v_CALCULATION_CNTR_2_port, Z => 
                           n1391);
   U4182 : ND2I port map( A => n4441, B => n3672, Z => n3708);
   U4183 : ND2I port map( A => v_CALCULATION_CNTR_2_port, B => n3671, Z => 
                           n3672);
   U4185 : ND2I port map( A => v_CALCULATION_CNTR_1_port, B => n1499, Z => 
                           n1498);
   U4193 : NR2I port map( A => RESET_I, B => n3954, Z => n1474);
   U4194 : ND2I port map( A => n3803, B => n4857, Z => n1483);
   U4196 : ND2I port map( A => v_CALCULATION_CNTR_2_port, B => n4601, Z => 
                           n2391);
   U4202 : ND2I port map( A => n4850, B => n4713, Z => n1454);
   KEXP0 : key_expansion port map( KEY_I(7) => KEY_I(7), KEY_I(6) => KEY_I(6), 
                           KEY_I(5) => KEY_I(5), KEY_I(4) => KEY_I(4), KEY_I(3)
                           => KEY_I(3), KEY_I(2) => KEY_I(2), KEY_I(1) => 
                           KEY_I(1), KEY_I(0) => KEY_I(0), VALID_KEY_I => 
                           VALID_KEY_I, CLK_I => CLK_I, RESET_I => RESET_I, 
                           CE_I => CE_I, DONE_O => KEY_READY_O, GET_KEY_I => 
                           GET_KEY, KEY_NUMB_I(5) => v_INV_KEY_NUMB_5_port, 
                           KEY_NUMB_I(4) => v_INV_KEY_NUMB_4_port, 
                           KEY_NUMB_I(3) => v_INV_KEY_NUMB_3_port, 
                           KEY_NUMB_I(2) => v_INV_KEY_NUMB_2_port, 
                           KEY_NUMB_I(1) => n4653, KEY_NUMB_I(0) => n4620, 
                           KEY_EXP_O(31) => v_KEY_COLUMN_31_port, KEY_EXP_O(30)
                           => v_KEY_COLUMN_30_port, KEY_EXP_O(29) => 
                           v_KEY_COLUMN_29_port, KEY_EXP_O(28) => 
                           v_KEY_COLUMN_28_port, KEY_EXP_O(27) => 
                           v_KEY_COLUMN_27_port, KEY_EXP_O(26) => 
                           v_KEY_COLUMN_26_port, KEY_EXP_O(25) => 
                           v_KEY_COLUMN_25_port, KEY_EXP_O(24) => 
                           v_KEY_COLUMN_24_port, KEY_EXP_O(23) => 
                           v_KEY_COLUMN_23_port, KEY_EXP_O(22) => 
                           v_KEY_COLUMN_22_port, KEY_EXP_O(21) => 
                           v_KEY_COLUMN_21_port, KEY_EXP_O(20) => 
                           v_KEY_COLUMN_20_port, KEY_EXP_O(19) => 
                           v_KEY_COLUMN_19_port, KEY_EXP_O(18) => 
                           v_KEY_COLUMN_18_port, KEY_EXP_O(17) => 
                           v_KEY_COLUMN_17_port, KEY_EXP_O(16) => 
                           v_KEY_COLUMN_16_port, KEY_EXP_O(15) => 
                           v_KEY_COLUMN_15_port, KEY_EXP_O(14) => 
                           v_KEY_COLUMN_14_port, KEY_EXP_O(13) => 
                           v_KEY_COLUMN_13_port, KEY_EXP_O(12) => 
                           v_KEY_COLUMN_12_port, KEY_EXP_O(11) => 
                           v_KEY_COLUMN_11_port, KEY_EXP_O(10) => 
                           v_KEY_COLUMN_10_port, KEY_EXP_O(9) => 
                           v_KEY_COLUMN_9_port, KEY_EXP_O(8) => 
                           v_KEY_COLUMN_8_port, KEY_EXP_O(7) => 
                           v_KEY_COLUMN_7_port, KEY_EXP_O(6) => 
                           v_KEY_COLUMN_6_port, KEY_EXP_O(5) => 
                           v_KEY_COLUMN_5_port, KEY_EXP_O(4) => 
                           v_KEY_COLUMN_4_port, KEY_EXP_O(3) => 
                           v_KEY_COLUMN_3_port, KEY_EXP_O(2) => 
                           v_KEY_COLUMN_2_port, KEY_EXP_O(1) => 
                           v_KEY_COLUMN_1_port, KEY_EXP_O(0) => 
                           v_KEY_COLUMN_0_port);
   U4205 : ND2I port map( A => n1467, B => n4462, Z => n4349);
   U4206 : NR2I port map( A => n103, B => n3939, Z => n4350);
   U4207 : NR2I port map( A => n4380, B => n103, Z => n4351);
   U4208 : ND2I port map( A => n4860, B => n4441, Z => n4352);
   U4209 : IVDA port map( A => n105, Y => n4353, Z => n4354);
   U4210 : AN2I port map( A => v_RAM_OUT0_20_port, B => n4365, Z => n4355);
   U4211 : AN2I port map( A => v_RAM_OUT0_4_port, B => n4363, Z => n4356);
   U4212 : AN2I port map( A => v_RAM_OUT0_28_port, B => n4362, Z => n4357);
   U4213 : ND3 port map( A => n4462, B => n1465, C => n3946, Z => n4358);
   U4214 : ND2I port map( A => n4378, B => n4404, Z => n4359);
   U4215 : ND2I port map( A => v_RAM_OUT0_12_port, B => n4378, Z => n4361);
   U4216 : EON1 port map( A => n4407, B => n1454, C => N2083, D => n1450, Z => 
                           n4309);
   U4217 : AN2I port map( A => v_RAM_OUT0_18_port, B => n4364, Z => n4369);
   U4218 : AN2I port map( A => v_RAM_OUT0_2_port, B => n4367, Z => n4370);
   U4219 : AN2I port map( A => v_RAM_OUT0_26_port, B => n4368, Z => n4371);
   U4220 : AN2I port map( A => v_RAM_OUT0_26_port, B => v_RAM_OUT0_28_port, Z 
                           => n4372);
   U4221 : AN2I port map( A => v_RAM_OUT0_2_port, B => v_RAM_OUT0_4_port, Z => 
                           n4373);
   U4222 : AN2I port map( A => v_RAM_OUT0_18_port, B => v_RAM_OUT0_20_port, Z 
                           => n4374);
   U4223 : ND2I port map( A => n3945, B => n1467, Z => n4375);
   U4224 : ND3 port map( A => n1465, B => n3946, C => n3945, Z => n4376);
   U4225 : NR3 port map( A => n4713, B => n3940, C => n4380, Z => n4377);
   U4226 : AN2I port map( A => v_RAM_OUT0_10_port, B => v_RAM_OUT0_12_port, Z 
                           => n4379);
   U4227 : ND3 port map( A => n4602, B => n4380, C => CE_I, Z => n4381);
   U4228 : NR4 port map( A => n4851, B => n4353, C => n1351, D => n1354, Z => 
                           n4382);
   U4229 : ND4 port map( A => n4860, B => n4354, C => n4856, D => n4850, Z => 
                           n4383);
   U4230 : AN3 port map( A => n1350, B => n4354, C => n1354, Z => n4386);
   U4231 : AN2I port map( A => n4366, B => n4859, Z => n4389);
   U4232 : NR3 port map( A => n4353, B => RESET_I, C => n4856, Z => n4496);
   U4233 : IVI port map( A => n4389, Z => n4706);
   U4234 : AO4 port map( A => n4754, B => n192_port, C => n4755, D => n4770, Z 
                           => n190);
   U4235 : AO4 port map( A => n4754, B => n4770, C => n4755, D => n192_port, Z 
                           => n188);
   U4236 : AO4 port map( A => n4748, B => n197, C => n199_port, D => n1003, Z 
                           => n1001);
   U4237 : AO4 port map( A => n197, B => n1003, C => n4748, D => n199_port, Z 
                           => n1004);
   U4238 : AO2 port map( A => n4360, B => n4975, C => n4702, D => n4969, Z => 
                           n2418);
   U4239 : AO4 port map( A => n4750, B => n4734, C => n4749, D => n661, Z => 
                           n1366);
   U4240 : AO4 port map( A => n4750, B => n661, C => n4749, D => n4734, Z => 
                           n1365);
   U4241 : AO4 port map( A => n1371, B => n197, C => n199_port, D => n4751, Z 
                           => n1370);
   U4242 : AO4 port map( A => n197, B => n4751, C => n1371, D => n199_port, Z 
                           => n1374);
   U4243 : AO4 port map( A => n196, B => n197, C => n4782, D => n199_port, Z =>
                           n195);
   U4244 : AO4 port map( A => n4782, B => n197, C => n196, D => n199_port, Z =>
                           n202_port);
   U4245 : IVI port map( A => n4386, Z => n4712);
   U4246 : EON1 port map( A => n4383, B => n1245, C => n4386, D => n4654, Z => 
                           n1243);
   U4247 : ENI port map( A => n1265, B => n1266, Z => n4654);
   U4248 : AO2 port map( A => n2995, B => n4355, C => n4374, D => n4948, Z => 
                           n3065);
   U4249 : AO2 port map( A => n3396, B => n4356, C => n4373, D => n5030, Z => 
                           n3467);
   U4250 : IVI port map( A => n2183, Z => n5040);
   U4251 : EO1 port map( A => n4876, B => n4357, C => n2503, D => n4705, Z => 
                           n2837);
   U4252 : EO1 port map( A => n4932, B => n4355, C => n2907, D => n4700, Z => 
                           n3241);
   U4253 : EON1 port map( A => n4918, B => n4700, C => n3089, D => n4355, Z => 
                           n3088);
   U4254 : AO2 port map( A => n4360, B => n4969, C => n2159, D => n4379, Z => 
                           n2252);
   U4255 : AO4 port map( A => n2211, B => n4361, C => n4359, D => n2212, Z => 
                           n2208);
   U4256 : AO4 port map( A => n4985, B => n4707, C => n2089_port, D => n4359, Z
                           => n2085_port);
   U4257 : EO1 port map( A => n5014, B => n4356, C => n3309, D => n4697, Z => 
                           n3643);
   U4258 : EON1 port map( A => n5000, B => n4697, C => n3491, D => n4356, Z => 
                           n3490);
   U4259 : AO2 port map( A => n4701, B => n4959, C => n4360, D => n4977, Z => 
                           n2417);
   U4260 : EO1 port map( A => n4360, B => n2190, C => n4361, D => n2191, Z => 
                           n2189);
   U4261 : AO2 port map( A => n2593, B => n4357, C => n4372, D => n4891, Z => 
                           n2660);
   U4262 : IVI port map( A => n2318, Z => n5041);
   U4263 : AO4 port map( A => n4361, B => n2133, C => n2199, D => n4707, Z => 
                           n2198);
   U4264 : AO7 port map( A => n4359, B => n2067, C => n4506, Z => n2197);
   U4265 : AO7 port map( A => n2874, B => n4371, C => n4884, Z => n2873);
   U4266 : AO7 port map( A => n3288, B => n4369, C => n4938, Z => n3287);
   U4267 : AO2 port map( A => n2048, B => n4360, C => n4379, D => n4977, Z => 
                           n2343);
   U4268 : AO7 port map( A => n3692, B => n4370, C => n5020, Z => n3691);
   U4269 : AO4 port map( A => n4889, B => n4704, C => n1958, D => n1959, Z => 
                           n1952);
   U4270 : EON1 port map( A => n4885, B => n4705, C => n2684, D => n4357, Z => 
                           n2683);
   U4271 : AO4 port map( A => n4949, B => n4698, C => n1689, D => n2957, Z => 
                           n3198);
   U4272 : AO4 port map( A => n4698, B => n2947, C => n4932, D => n2957, Z => 
                           n3087);
   U4273 : AO4 port map( A => n4918, B => n4698, C => n2957, D => n3095, Z => 
                           n3091);
   U4274 : AO4 port map( A => n4700, B => n3093, C => n3094, D => n4682, Z => 
                           n3092);
   U4275 : AO4 port map( A => n2372, B => n4359, C => n4978, D => n4361, Z => 
                           n2405);
   U4276 : EON1 port map( A => n4361, B => n2166, C => n2056, D => n4702, Z => 
                           n2163);
   U4277 : AO4 port map( A => n5031, B => n4695, C => n2455, D => n3359, Z => 
                           n3599);
   U4278 : AO4 port map( A => n4695, B => n3349, C => n5014, D => n3359, Z => 
                           n3489);
   U4279 : AO4 port map( A => n5000, B => n4695, C => n3359, D => n3497, Z => 
                           n3493);
   U4280 : AO4 port map( A => n4697, B => n3495, C => n3496, D => n4678, Z => 
                           n3494);
   U4281 : AO2 port map( A => n5042, B => n2796, C => n4399, D => n2797, Z => 
                           n2795);
   U4282 : AO3 port map( A => n2755, B => n4705, C => n2660, D => n2801, Z => 
                           n2796);
   U4283 : AO3 port map( A => n4704, B => n2654, C => n2798, D => n2799, Z => 
                           n2797);
   U4284 : AO2 port map( A => n4703, B => n2802, C => n4887, D => n4372, Z => 
                           n2801);
   U4285 : AO2 port map( A => n5037, B => n3214, C => n4402, D => n3215, Z => 
                           n3213);
   U4286 : AO3 port map( A => n3159, B => n4700, C => n3065, D => n3219, Z => 
                           n3214);
   U4287 : AO3 port map( A => n4698, B => n3058, C => n3216, D => n3217, Z => 
                           n3215);
   U4288 : AO2 port map( A => n4699, B => n3220, C => n4928, D => n4374, Z => 
                           n3219);
   U4289 : AO2 port map( A => n5044, B => n3615, C => n4400, D => n3616, Z => 
                           n3614);
   U4290 : AO3 port map( A => n3560, B => n4697, C => n3467, D => n3620, Z => 
                           n3615);
   U4291 : AO3 port map( A => n4695, B => n3460, C => n3617, D => n3618, Z => 
                           n3616);
   U4292 : AO2 port map( A => n4696, B => n3621, C => n5010, D => n4373, Z => 
                           n3620);
   U4293 : AO2 port map( A => n4702, B => n2192, C => n4983, D => n4379, Z => 
                           n2188);
   U4294 : AO4 port map( A => n4704, B => n2649, C => n4882, D => n1959, Z => 
                           n2847);
   U4295 : AO2 port map( A => n2755, B => n4703, C => n2707, D => n4372, Z => 
                           n2754);
   U4296 : AO4 port map( A => n4698, B => n3053, C => n4954, D => n2957, Z => 
                           n3251);
   U4297 : AO2 port map( A => n3159, B => n4699, C => n3112, D => n4374, Z => 
                           n3158);
   U4298 : AO4 port map( A => n4707, B => n2190, C => n4995, D => n4359, Z => 
                           n2360);
   U4299 : AO4 port map( A => n4695, B => n3455, C => n5036, D => n3359, Z => 
                           n3653);
   U4300 : AO2 port map( A => n3560, B => n4696, C => n3513, D => n4373, Z => 
                           n3559);
   U4301 : IVI port map( A => n4372, Z => n4704);
   U4302 : IVI port map( A => n4374, Z => n4698);
   U4303 : IVI port map( A => n4369, Z => n4700);
   U4304 : AO4 port map( A => n4704, B => n2542, C => n4876, D => n1959, Z => 
                           n2682);
   U4305 : AO4 port map( A => n4885, B => n4704, C => n1959, D => n2690, Z => 
                           n2686);
   U4306 : AO4 port map( A => n4705, B => n2688, C => n2689, D => n4687, Z => 
                           n2687);
   U4307 : AO4 port map( A => n4361, B => n4958, C => n2179, D => n4690, Z => 
                           n2342);
   U4308 : AO4 port map( A => n4985, B => n4690, C => n2293, D => n4361, Z => 
                           n2359);
   U4309 : AO4 port map( A => n4985, B => n4690, C => n5069, D => n4361, Z => 
                           n2300);
   U4310 : IVI port map( A => n4373, Z => n4695);
   U4311 : AO2 port map( A => n4357, B => n4897, C => n4703, D => n2761, Z => 
                           n2799);
   U4312 : AO2 port map( A => n4355, B => n5066, C => n4699, D => n3165, Z => 
                           n3217);
   U4313 : AO2 port map( A => n4356, B => n5071, C => n4696, D => n3566, Z => 
                           n3618);
   U4314 : AO4 port map( A => n4705, B => n2533, C => n2652, D => n4687, Z => 
                           n2805);
   U4315 : AO4 port map( A => n4700, B => n2939, C => n3056, D => n4682, Z => 
                           n3224);
   U4316 : AO4 port map( A => n2158, B => n4707, C => n4980, D => n4359, Z => 
                           n2346);
   U4317 : EON1 port map( A => n4995, B => n4690, C => n2140, D => n4701, Z => 
                           n2345);
   U4318 : AO4 port map( A => n4697, B => n3341, C => n3458, D => n4678, Z => 
                           n3625);
   U4319 : AO2 port map( A => n4900, B => n5062, C => n5061, D => n2678, Z => 
                           n2856);
   U4320 : AO2 port map( A => n4941, B => n5054, C => n5053, D => n3083, Z => 
                           n3260);
   U4321 : AO2 port map( A => n5023, B => n5048, C => n5047, D => n3485, Z => 
                           n3662);
   U4322 : AO4 port map( A => n4872, B => n4705, C => n2756, D => n4687, Z => 
                           n2848);
   U4323 : AO2 port map( A => n2756, B => n4357, C => n4883, D => n4371, Z => 
                           n2753);
   U4324 : AO4 port map( A => n4944, B => n4700, C => n3160, D => n4682, Z => 
                           n3252);
   U4325 : AO2 port map( A => n3160, B => n4355, C => n5065, D => n4369, Z => 
                           n3157);
   U4326 : AO4 port map( A => n5026, B => n4697, C => n3561, D => n4678, Z => 
                           n3654);
   U4327 : AO2 port map( A => n3561, B => n4356, C => n5070, D => n4370, Z => 
                           n3558);
   U4328 : AO4 port map( A => n4747, B => n998, C => n4746, D => n4765, Z => 
                           n996);
   U4329 : AO4 port map( A => n4747, B => n4765, C => n4746, D => n998, Z => 
                           n994);
   U4330 : AO4 port map( A => n4712, B => n760, C => n4383, D => n761, Z => 
                           n759);
   U4331 : AO4 port map( A => n4712, B => n503, C => n4383, D => n504, Z => 
                           n502);
   U4332 : AO4 port map( A => n4712, B => n934, C => n4383, D => n935, Z => 
                           n933);
   U4333 : AO4 port map( A => n4712, B => n330, C => n4383, D => n331, Z => 
                           n329);
   U4334 : AO4 port map( A => n4712, B => n1168, C => n4383, D => n1169, Z => 
                           n1167);
   U4335 : AO4 port map( A => n4712, B => n839, C => n4383, D => n840, Z => 
                           n838);
   U4336 : AO4 port map( A => n4712, B => n528, C => n4383, D => n529, Z => 
                           n527);
   U4337 : AO4 port map( A => n4712, B => n567, C => n4383, D => n568, Z => 
                           n566);
   U4338 : AO4 port map( A => n4712, B => n113, C => n4383, D => n115, Z => 
                           n111);
   U4339 : AO4 port map( A => n4712, B => n797, C => n4383, D => n798, Z => 
                           n796);
   U4340 : AO4 port map( A => n4712, B => n892, C => n4383, D => n893, Z => 
                           n891);
   U4341 : AO4 port map( A => n4712, B => n264, C => n4383, D => n265, Z => 
                           n263);
   U4342 : AO4 port map( A => n4712, B => n1040, C => n4383, D => n1041, Z => 
                           n1039);
   U4343 : AO4 port map( A => n4712, B => n706, C => n4383, D => n707, Z => 
                           n705);
   U4344 : AO4 port map( A => n4712, B => n396, C => n4383, D => n397, Z => 
                           n395);
   U4345 : AO4 port map( A => n4712, B => n668, C => n4383, D => n669, Z => 
                           n667);
   U4346 : AO4 port map( A => n4712, B => n371, C => n4383, D => n372, Z => 
                           n370);
   U4347 : AO4 port map( A => n4712, B => n625, C => n4383, D => n626, Z => 
                           n624);
   U4348 : AO3 port map( A => n4361, B => n4978, C => n2421, D => n2110, Z => 
                           n2410);
   U4349 : AO2 port map( A => n4910, B => n2414, C => n4909, D => n2415, Z => 
                           n2413);
   U4350 : AO3 port map( A => n4361, B => n2144, C => n2087_port, D => n2418, Z
                           => n2414);
   U4351 : EO1 port map( A => n4702, B => n2098, C => n2144, D => n4707, Z => 
                           n2416);
   U4352 : AO3 port map( A => n4938, B => n2936, C => n2981, D => n2982, Z => 
                           n2979);
   U4353 : EO1 port map( A => n2993, B => n5057, C => n2995, D => n2940, Z => 
                           n2981);
   U4354 : EON1 port map( A => n2988, B => n2989, C => n2990, D => n2926, Z => 
                           n2984);
   U4355 : IVDA port map( A => n3708, Y => n4366, Z => n4673);
   U4356 : AO3 port map( A => n4905, B => n4569, C => n2316, D => n2317, Z => 
                           n1549);
   U4357 : AO3 port map( A => n4986, B => n2318, C => n2327, D => n2328, Z => 
                           n2316);
   U4358 : EON1 port map( A => n2331, B => n4690, C => n2067, D => n4701, Z => 
                           n2381);
   U4359 : AO3 port map( A => n4884, B => n2530, C => n2578, D => n2579, Z => 
                           n2577);
   U4360 : EO1 port map( A => n2591, B => n5060, C => n2593, D => n2534, Z => 
                           n2578);
   U4361 : AO3 port map( A => n5020, B => n3338, C => n3382, D => n3383, Z => 
                           n3380);
   U4362 : EO1 port map( A => n3394, B => n5051, C => n3396, D => n3342, Z => 
                           n3382);
   U4363 : NR4 port map( A => n3049, B => n4919, C => n3051, D => n3052, Z => 
                           n3048);
   U4364 : EON1 port map( A => n2947, B => n3055, C => n2938, D => n3056, Z => 
                           n3051);
   U4365 : AO4 port map( A => n2988, B => n3053, C => n4954, D => n2936, Z => 
                           n3052);
   U4366 : AO3 port map( A => n3060, B => n2923, C => n3061, D => n4409, Z => 
                           n3049);
   U4367 : NR4 port map( A => n3451, B => n5001, C => n3453, D => n3454, Z => 
                           n3450);
   U4368 : EON1 port map( A => n3349, B => n3457, C => n3340, D => n3458, Z => 
                           n3453);
   U4369 : AO4 port map( A => n3389, B => n3455, C => n5036, D => n3338, Z => 
                           n3454);
   U4370 : AO3 port map( A => n3462, B => n3325, C => n3463, D => n4408, Z => 
                           n3451);
   U4371 : ND4 port map( A => n2878, B => n2879, C => n2880, D => n2881, Z => 
                           n1982);
   U4372 : AO2 port map( A => n5061, B => n2618, C => n2522, D => n2552, Z => 
                           n2880);
   U4373 : AO2 port map( A => n2531, B => n4880, C => n5060, D => n4913, Z => 
                           n2878);
   U4374 : ND4 port map( A => n3289, B => n3290, C => n3291, D => n3292, Z => 
                           n1705);
   U4375 : AO2 port map( A => n5053, B => n3020, C => n2926, D => n2955, Z => 
                           n3291);
   U4376 : AO2 port map( A => n2938, B => n4933, C => n5057, D => n4937, Z => 
                           n3289);
   U4377 : ND4 port map( A => n3693, B => n3694, C => n3695, D => n3696, Z => 
                           n2469);
   U4378 : AO2 port map( A => n5047, B => n3421, C => n3328, D => n3357, Z => 
                           n3695);
   U4379 : AO2 port map( A => n3340, B => n5015, C => n5051, D => n5019, Z => 
                           n3693);
   U4380 : AO2 port map( A => n4360, B => n2203, C => n2234, D => n4702, Z => 
                           n2312);
   U4381 : EON1 port map( A => n2585, B => n2586, C => n2587, D => n2522, Z => 
                           n2581);
   U4382 : AO2 port map( A => n2525, B => n4511, C => n2527, D => n2528, Z => 
                           n2520);
   U4383 : AO2 port map( A => n2930, B => n4512, C => n2932, D => n2933, Z => 
                           n2924);
   U4384 : AO4 port map( A => n4707, B => n4974, C => n2150, D => n4690, Z => 
                           n2147);
   U4385 : EON1 port map( A => n3389, B => n3390, C => n3391, D => n3328, Z => 
                           n3385);
   U4386 : AO2 port map( A => n3332, B => n4513, C => n3334, D => n3335, Z => 
                           n3326);
   U4387 : AO2 port map( A => n4503, B => n2832, C => n4399, D => n2833, Z => 
                           n2831);
   U4388 : AO7 port map( A => n4687, B => n2738, C => n2834, Z => n2833);
   U4389 : AO3 port map( A => n4704, B => n2540, C => n2836, D => n2837, Z => 
                           n2832);
   U4390 : AO2 port map( A => n4504, B => n3236, C => n4402, D => n3237, Z => 
                           n3235);
   U4391 : AO7 port map( A => n4682, B => n3142, C => n3238, Z => n3237);
   U4392 : AO3 port map( A => n4698, B => n1722, C => n3240, D => n3241, Z => 
                           n3236);
   U4393 : EO1 port map( A => n3239, B => n1722, C => n3011, D => n2957, Z => 
                           n3238);
   U4394 : AO3 port map( A => n3084, B => n4685, C => n3085, D => n3086, Z => 
                           n3044);
   U4395 : AO7 port map( A => n3091, B => n3092, C => n5037, Z => n3085);
   U4396 : AO7 port map( A => n3087, B => n3088, C => n5038, Z => n3086);
   U4397 : AO4 port map( A => n2298, B => n4691, C => n2299, D => n1897, Z => 
                           n2297);
   U4398 : AO6 port map( A => n2084_port, B => n4379, C => n2302, Z => n2298);
   U4399 : AO4 port map( A => n4997, B => n4690, C => n2304, D => n2305, Z => 
                           n2302);
   U4400 : AO2 port map( A => n5069, B => n2292, C => n2293, D => n2054, Z => 
                           n2286);
   U4401 : AO4 port map( A => n2201, B => n2074, C => n2202, D => n1912, Z => 
                           n2195);
   U4402 : AO4 port map( A => n4359, B => n2044, C => n2206, D => n4361, Z => 
                           n2204);
   U4403 : AO4 port map( A => n2138, B => n4691, C => n2139, D => n1897, Z => 
                           n2137);
   U4404 : AO4 port map( A => n2082, B => n1897, C => n2083_port, D => n4691, Z
                           => n2070);
   U4405 : AO7 port map( A => n4378, B => n4981, C => n4690, Z => n2090);
   U4406 : AO2 port map( A => n4505, B => n3638, C => n4400, D => n3639, Z => 
                           n3637);
   U4407 : AO7 port map( A => n4678, B => n3543, C => n3640, Z => n3639);
   U4408 : AO3 port map( A => n4695, B => n2486, C => n3642, D => n3643, Z => 
                           n3638);
   U4409 : EO1 port map( A => n3641, B => n2486, C => n3412, D => n3359, Z => 
                           n3640);
   U4410 : AO3 port map( A => n3486, B => n4681, C => n3487, D => n3488, Z => 
                           n3446);
   U4411 : AO7 port map( A => n3493, B => n3494, C => n5044, Z => n3487);
   U4412 : AO7 port map( A => n3489, B => n3490, C => n5045, Z => n3488);
   U4413 : AO4 port map( A => n4707, B => n2120, C => n2210, D => n4359, Z => 
                           n2301);
   U4414 : AO7 port map( A => n4669, B => n4706, C => n1923, Z => n1934);
   U4415 : AO7 port map( A => v_KEY_COLUMN_29_port, B => n4706, C => n1923, Z 
                           => n1930);
   U4416 : AO7 port map( A => n4671, B => n4706, C => n1923, Z => n1922);
   U4417 : AO7 port map( A => v_KEY_COLUMN_0_port, B => n4706, C => n2426, Z =>
                           n2466);
   U4418 : AO7 port map( A => v_KEY_COLUMN_2_port, B => n4706, C => n2426, Z =>
                           n2440);
   U4419 : AO7 port map( A => n4667, B => n1527, C => n2495, Z => n2865);
   U4420 : AO7 port map( A => v_KEY_COLUMN_26_port, B => n1527, C => n2495, Z 
                           => n2790);
   U4421 : AO7 port map( A => n4664, B => n1527, C => n2897, Z => n3103);
   U4422 : AO7 port map( A => n4665, B => n1527, C => n2897, Z => n2974);
   U4423 : AO7 port map( A => v_KEY_COLUMN_16_port, B => n1609, C => n1650, Z 
                           => n1701);
   U4424 : AO7 port map( A => v_KEY_COLUMN_18_port, B => n1609, C => n1650, Z 
                           => n1674);
   U4425 : AO7 port map( A => v_KEY_COLUMN_1_port, B => n1609, C => n1759, Z =>
                           n1779);
   U4426 : AO7 port map( A => n4655, B => n1609, C => n1759, Z => n1766);
   U4427 : AO2 port map( A => n3053, B => n2926, C => n3058, D => n5053, Z => 
                           n3057);
   U4428 : AO2 port map( A => n3455, B => n3328, C => n3460, D => n5047, Z => 
                           n3459);
   U4429 : AO4 port map( A => n4359, B => n2154, C => n4707, D => n2382, Z => 
                           n2205);
   U4430 : AO6 port map( A => n2528, B => n2583, C => n4705, Z => n2777);
   U4431 : AO4 port map( A => n4687, B => n2593, C => n2601, D => n1959, Z => 
                           n2776);
   U4432 : AO6 port map( A => n2933, B => n2986, C => n4700, Z => n3181);
   U4433 : AO4 port map( A => n4682, B => n2995, C => n3003, D => n2957, Z => 
                           n3180);
   U4434 : AO6 port map( A => n2167, B => n2212, C => n4361, Z => n2379);
   U4435 : AO4 port map( A => n4707, B => n1907, C => n4985, D => n4359, Z => 
                           n2378);
   U4436 : AO6 port map( A => n3335, B => n3387, C => n4697, Z => n3582);
   U4437 : AO4 port map( A => n4678, B => n3396, C => n3404, D => n3359, Z => 
                           n3581);
   U4438 : AO3 port map( A => n2532, B => n2530, C => n2778, D => n2779, Z => 
                           n2769);
   U4439 : AO2 port map( A => n5060, B => n2785, C => n4878, D => n2531, Z => 
                           n2778);
   U4440 : AO3 port map( A => n3182, B => n2936, C => n3183, D => n3184, Z => 
                           n3173);
   U4441 : AO2 port map( A => n5057, B => n3190, C => n4940, D => n2938, Z => 
                           n3183);
   U4442 : AO4 port map( A => n4682, B => n2965, C => n2957, D => n3039, Z => 
                           n3037);
   U4443 : NR3 port map( A => n4700, B => n4935, C => n4926, Z => n3038);
   U4444 : AO3 port map( A => n3583, B => n3338, C => n3584, D => n3585, Z => 
                           n3574);
   U4445 : AO2 port map( A => n5051, B => n3591, C => n5022, D => n3340, Z => 
                           n3584);
   U4446 : NR4 port map( A => n2645, B => n4877, C => n2647, D => n2648, Z => 
                           n2644);
   U4447 : EON1 port map( A => n2542, B => n2651, C => n2531, D => n2652, Z => 
                           n2647);
   U4448 : AO4 port map( A => n2585, B => n2649, C => n4882, D => n2530, Z => 
                           n2648);
   U4449 : AO3 port map( A => n2655, B => n2519, C => n2656, D => n4410, Z => 
                           n2645);
   U4450 : ND4 port map( A => n2817, B => n2818, C => n2819, D => n2820, Z => 
                           n1944);
   U4451 : AO2 port map( A => n2522, B => n2822, C => n5060, D => n2529, Z => 
                           n2818);
   U4452 : AO2 port map( A => n2707, B => n5062, C => n5061, D => n2621, Z => 
                           n2819);
   U4453 : AO2 port map( A => n2531, B => n2821, C => n2527, D => n4686, Z => 
                           n2820);
   U4454 : ND4 port map( A => n3203, B => n3204, C => n3205, D => n3206, Z => 
                           n1679);
   U4455 : AO2 port map( A => n2926, B => n3208, C => n5057, D => n2935, Z => 
                           n3204);
   U4456 : AO2 port map( A => n3112, B => n5054, C => n5053, D => n3024, Z => 
                           n3205);
   U4457 : AO2 port map( A => n2938, B => n3207, C => n2932, D => n4683, Z => 
                           n3206);
   U4458 : ND4 port map( A => n3604, B => n3605, C => n3606, D => n3607, Z => 
                           n2445);
   U4459 : AO2 port map( A => n3328, B => n3609, C => n5051, D => n3337, Z => 
                           n3605);
   U4460 : AO2 port map( A => n3513, B => n5048, C => n5047, D => n3425, Z => 
                           n3606);
   U4461 : AO2 port map( A => n3340, B => n3608, C => n3334, D => n4679, Z => 
                           n3607);
   U4462 : AO7 port map( A => n4890, B => n4881, C => n4371, Z => n2798);
   U4463 : AO7 port map( A => n4365, B => n3095, C => n4700, Z => n3239);
   U4464 : AO7 port map( A => n4936, B => n4942, C => n4369, Z => n3216);
   U4465 : AO6 port map( A => n2283, B => n4378, C => n4702, Z => n2304);
   U4466 : AO7 port map( A => n4363, B => n3497, C => n4697, Z => n3641);
   U4467 : AO7 port map( A => n5018, B => n5024, C => n4370, Z => n3617);
   U4468 : EO1 port map( A => n2835, B => n2540, C => n2608, D => n1959, Z => 
                           n2834);
   U4469 : AO7 port map( A => n4362, B => n2690, C => n4705, Z => n2835);
   U4470 : AO2 port map( A => n2522, B => n2523, C => n5059, D => n4895, Z => 
                           n2521);
   U4471 : AO4 port map( A => n2968, B => n4700, C => n4946, D => n2957, Z => 
                           n3096);
   U4472 : AO6 port map( A => n2957, B => n3002, C => n3003, Z => n3000);
   U4473 : AO2 port map( A => n2926, B => n2927, C => n5056, D => n4939, Z => 
                           n2925);
   U4474 : AO4 port map( A => n4956, B => n1912, C => n1916, D => n4691, Z => 
                           n1910);
   U4475 : AO4 port map( A => n4707, B => n1913, C => n2046, D => n4359, Z => 
                           n2361);
   U4476 : EON1 port map( A => n4359, B => n2154, C => n2166, D => n4379, Z => 
                           n2387);
   U4477 : AO4 port map( A => n1901, B => n2281, C => n4361, D => n2060, Z => 
                           n2349);
   U4478 : AO4 port map( A => n4690, B => n2144, C => n2145, D => n4361, Z => 
                           n2141);
   U4479 : AO7 port map( A => n2113, B => n4690, C => n2165, Z => n2164);
   U4480 : AO4 port map( A => n2128, B => n4707, C => n4690, D => n4996, Z => 
                           n2127);
   U4481 : AO4 port map( A => n3370, B => n4697, C => n5028, D => n3359, Z => 
                           n3498);
   U4482 : AO2 port map( A => n3328, B => n3329, C => n5050, D => n5021, Z => 
                           n3327);
   U4483 : AO2 port map( A => n4984, B => n5041, C => n5040, D => n1907, Z => 
                           n2396);
   U4484 : AO2 port map( A => n5059, B => n2861, C => n2527, D => n2850, Z => 
                           n2857);
   U4485 : AO2 port map( A => n5063, B => n4880, C => n5059, D => n2528, Z => 
                           n2817);
   U4486 : AO2 port map( A => n5056, B => n3265, C => n2932, D => n3254, Z => 
                           n3261);
   U4487 : AO2 port map( A => n5055, B => n4933, C => n5056, D => n2933, Z => 
                           n3203);
   U4488 : AO2 port map( A => n2926, B => n2964, C => n1689, D => n2938, Z => 
                           n2997);
   U4489 : AO3 port map( A => n4359, B => n2380, C => n2420, D => n1878, Z => 
                           n2419);
   U4490 : AO2 port map( A => n5050, B => n3667, C => n3334, D => n3656, Z => 
                           n3663);
   U4491 : AO2 port map( A => n5049, B => n5015, C => n5050, D => n3335, Z => 
                           n3604);
   U4492 : AO4 port map( A => n4874, B => n4689, C => n1985, D => n4688, Z => 
                           n1983);
   U4493 : AO6 port map( A => n1978, B => n1986, C => n1987, Z => n1985);
   U4494 : AO4 port map( A => n4705, B => n1988, C => n4885, D => n4687, Z => 
                           n1987);
   U4495 : AO4 port map( A => n2845, B => n4688, C => n2846, D => n4689, Z => 
                           n2844);
   U4496 : AO6 port map( A => n2529, B => n2714, C => n4705, Z => n2852);
   U4497 : AO3 port map( A => n2762, B => n2530, C => n2763, D => n2764, Z => 
                           n2748);
   U4498 : AO2 port map( A => n2767, B => n5061, C => n2531, D => n2768, Z => 
                           n2763);
   U4499 : AO2 port map( A => n5059, B => n2765, C => n4888, D => n2527, Z => 
                           n2764);
   U4500 : AO3 port map( A => n2679, B => n4688, C => n2680, D => n2681, Z => 
                           n2640);
   U4501 : AO7 port map( A => n2686, B => n2687, C => n5042, Z => n2680);
   U4502 : AO7 port map( A => n2682, B => n2683, C => n5043, Z => n2681);
   U4503 : AO4 port map( A => n2501, B => n4689, C => n2502, D => n4688, Z => 
                           n2500);
   U4504 : AO6 port map( A => n2503, B => n4362, C => n2505, Z => n2502);
   U4505 : AO6 port map( A => n4703, B => n2509, C => n2510, Z => n2501);
   U4506 : AO4 port map( A => n4896, B => n4687, C => n2507, D => n4705, Z => 
                           n2505);
   U4507 : AO4 port map( A => n4924, B => n4684, C => n3282, D => n4685, Z => 
                           n3281);
   U4508 : AO6 port map( A => n1712, B => n1710, C => n3283, Z => n3282);
   U4509 : AO4 port map( A => n4700, B => n1713, C => n4918, D => n4682, Z => 
                           n3283);
   U4510 : AO4 port map( A => n3249, B => n4685, C => n3250, D => n4684, Z => 
                           n3248);
   U4511 : AO6 port map( A => n2935, B => n3118, C => n4700, Z => n3256);
   U4512 : AO3 port map( A => n3166, B => n2936, C => n3167, D => n3168, Z => 
                           n3152);
   U4513 : AO2 port map( A => n3171, B => n5053, C => n2938, D => n3172, Z => 
                           n3167);
   U4514 : AO2 port map( A => n5056, B => n3169, C => n4929, D => n2932, Z => 
                           n3168);
   U4515 : AO4 port map( A => n2903, B => n4684, C => n2905, D => n4685, Z => 
                           n2902);
   U4516 : AO6 port map( A => n2907, B => n4365, C => n2908, Z => n2905);
   U4517 : AO6 port map( A => n4699, B => n2913, C => n2914, Z => n2903);
   U4518 : AO4 port map( A => n4934, B => n4682, C => n2911, D => n4700, Z => 
                           n2908);
   U4519 : AO4 port map( A => n2357, B => n4691, C => n2358, D => n1897, Z => 
                           n2356);
   U4520 : NR3 port map( A => n4361, B => n4964, C => n4991, Z => n2362);
   U4521 : AO2 port map( A => n4989, B => n2065, C => n4973, D => n5041, Z => 
                           n2285);
   U4522 : AO2 port map( A => n2054, B => n2133, C => n2278, D => n2279, Z => 
                           n2272);
   U4523 : AO6 port map( A => n4379, B => n4994, C => n4516, Z => n2278);
   U4524 : AO3 port map( A => n2155, B => n4516, C => n2156, D => n2157, Z => 
                           n2136);
   U4525 : AO2 port map( A => n2160, B => n5039, C => n2065, D => n2162, Z => 
                           n2156);
   U4526 : AO2 port map( A => n2158, B => n5040, C => n2159, D => n5041, Z => 
                           n2157);
   U4527 : AO4 port map( A => n5006, B => n4680, C => n3686, D => n4681, Z => 
                           n3685);
   U4528 : AO6 port map( A => n2476, B => n2474, C => n3687, Z => n3686);
   U4529 : AO4 port map( A => n4697, B => n2477, C => n5000, D => n4678, Z => 
                           n3687);
   U4530 : AO4 port map( A => n3651, B => n4681, C => n3652, D => n4680, Z => 
                           n3650);
   U4531 : AO6 port map( A => n3337, B => n3519, C => n4697, Z => n3658);
   U4532 : AO3 port map( A => n3567, B => n3338, C => n3568, D => n3569, Z => 
                           n3553);
   U4533 : AO2 port map( A => n3572, B => n5047, C => n3340, D => n3573, Z => 
                           n3568);
   U4534 : AO2 port map( A => n5050, B => n3570, C => n5011, D => n3334, Z => 
                           n3569);
   U4535 : AO4 port map( A => n3305, B => n4680, C => n3307, D => n4681, Z => 
                           n3304);
   U4536 : AO6 port map( A => n3309, B => n4363, C => n3310, Z => n3307);
   U4537 : AO6 port map( A => n4696, B => n3315, C => n3316, Z => n3305);
   U4538 : AO4 port map( A => n5016, B => n4678, C => n3313, D => n4697, Z => 
                           n3310);
   U4539 : AO3 port map( A => n4687, B => n2619, C => n2872, D => n2873, Z => 
                           n2871);
   U4540 : AO3 port map( A => n4682, B => n3022, C => n3286, D => n3287, Z => 
                           n3285);
   U4541 : AO3 port map( A => n4678, B => n3423, C => n3690, D => n3691, Z => 
                           n3689);
   U4542 : AO3 port map( A => n2793, B => n2544, C => n2794, D => n2795, Z => 
                           n2792);
   U4543 : AO7 port map( A => n2804, B => n2805, C => n4503, Z => n2794);
   U4544 : AO3 port map( A => n3211, B => n2949, C => n3212, D => n3213, Z => 
                           n3210);
   U4545 : AO7 port map( A => n3223, B => n3224, C => n4504, Z => n3212);
   U4546 : AO3 port map( A => n2334, B => n1912, C => n2335, D => n2336, Z => 
                           n2333);
   U4547 : AO7 port map( A => n2345, B => n2346, C => n4909, Z => n2335);
   U4548 : AO3 port map( A => n3612, B => n3351, C => n3613, D => n3614, Z => 
                           n3611);
   U4549 : AO7 port map( A => n3624, B => n3625, C => n4505, Z => n3613);
   U4550 : AO2 port map( A => n2331, B => n4701, C => n4360, D => n2093, Z => 
                           n2330);
   U4551 : AO2 port map( A => n4702, B => n1907, C => n4973, D => n4379, Z => 
                           n2329);
   U4552 : AO2 port map( A => n4503, B => n2751, C => n4399, D => n2752, Z => 
                           n2750);
   U4553 : AO3 port map( A => n1959, B => n2540, C => n2757, D => n2758, Z => 
                           n2751);
   U4554 : AO2 port map( A => n4504, B => n3155, C => n4402, D => n3156, Z => 
                           n3154);
   U4555 : AO3 port map( A => n2957, B => n1722, C => n3161, D => n3162, Z => 
                           n3155);
   U4556 : AO2 port map( A => n4702, B => n4996, C => n4379, D => n4967, Z => 
                           n2096);
   U4557 : AO2 port map( A => n4701, B => n2098, C => n4360, D => n1900, Z => 
                           n2097);
   U4558 : AO2 port map( A => n4505, B => n3556, C => n4400, D => n3557, Z => 
                           n3555);
   U4559 : AO3 port map( A => n3359, B => n2486, C => n3562, D => n3563, Z => 
                           n3556);
   U4560 : AO2 port map( A => n2649, B => n2522, C => n2654, D => n5061, Z => 
                           n2653);
   U4561 : ND3 port map( A => n1688, B => n4365, C => n4683, Z => n2992);
   U4562 : IVI port map( A => n4371, Z => n4705);
   U4563 : IVI port map( A => n4370, Z => n4697);
   U4564 : AO4 port map( A => n4872, B => n4705, C => n4883, D => n4687, Z => 
                           n2773);
   U4565 : AO4 port map( A => n4944, B => n4700, C => n5065, D => n4682, Z => 
                           n3177);
   U4566 : AO4 port map( A => n5026, B => n4697, C => n5070, D => n4678, Z => 
                           n3578);
   U4567 : AO4 port map( A => n4687, B => n2562, C => n1959, D => n2635, Z => 
                           n2633);
   U4568 : NR3 port map( A => n4705, B => n4912, C => n4901, Z => n2634);
   U4569 : AO3 port map( A => n4690, B => n2075, C => n2076, D => n2077, Z => 
                           n2073);
   U4570 : AO7 port map( A => n4955, B => n5069, C => n4379, Z => n2076);
   U4571 : AO4 port map( A => n4678, B => n3367, C => n3359, D => n3440, Z => 
                           n3438);
   U4572 : NR3 port map( A => n4697, B => n5017, C => n5008, Z => n3439);
   U4573 : IVDA port map( A => n2043, Y => n4360, Z => n4690);
   U4574 : IVDA port map( A => n1513, Y => n4515, Z => n4674);
   U4575 : IVDA port map( A => n1520, Y => n4452, Z => n4676);
   U4576 : IVDA port map( A => n1521, Y => n4564, Z => n4675);
   U4577 : ND3 port map( A => n4863, B => n4384, C => n2019, Z => n1562);
   U4578 : AO6 port map( A => n2093, B => n2167, C => n4707, Z => n2340);
   U4579 : AO7 port map( A => n4997, B => n4990, C => n4379, Z => n2311);
   U4580 : AO4 port map( A => n2853, B => n1959, C => n4704, D => n2854, Z => 
                           n2851);
   U4581 : AO2 port map( A => n2591, B => n4357, C => n4371, D => n2590, Z => 
                           n2758);
   U4582 : AO2 port map( A => n2719, B => n4362, C => n4914, D => n4368, Z => 
                           n2718);
   U4583 : AO4 port map( A => n2565, B => n4705, C => n4915, D => n1959, Z => 
                           n2691);
   U4584 : AO6 port map( A => n1959, B => n2600, C => n2601, Z => n2598);
   U4585 : AO4 port map( A => n3257, B => n2957, C => n4698, D => n3258, Z => 
                           n3255);
   U4586 : AO2 port map( A => n2993, B => n4355, C => n4369, D => n1688, Z => 
                           n3162);
   U4587 : AO2 port map( A => n3123, B => n4365, C => n4925, D => n4364, Z => 
                           n3122);
   U4588 : AO2 port map( A => n4701, B => n2239, C => n2128, D => n4379, Z => 
                           n2238);
   U4589 : AO4 port map( A => n3659, B => n3359, C => n4695, D => n3660, Z => 
                           n3657);
   U4590 : AO2 port map( A => n3394, B => n4356, C => n4370, D => n2454, Z => 
                           n3563);
   U4591 : AO2 port map( A => n3524, B => n4363, C => n5007, D => n4367, Z => 
                           n3523);
   U4592 : AO6 port map( A => n3359, B => n3403, C => n3404, Z => n3401);
   U4593 : AO2 port map( A => n4899, B => n5063, C => n5061, D => n2808, Z => 
                           n2891);
   U4594 : AO2 port map( A => n2859, B => n2531, C => n2522, D => n2860, Z => 
                           n2858);
   U4595 : AO2 port map( A => n2522, B => n2561, C => n1958, D => n2531, Z => 
                           n2595);
   U4596 : AO2 port map( A => n4943, B => n5055, C => n5053, D => n3227, Z => 
                           n3275);
   U4597 : AO2 port map( A => n3263, B => n2938, C => n2926, D => n3264, Z => 
                           n3262);
   U4598 : AO4 port map( A => n4359, B => n2182, C => n4361, D => n1913, Z => 
                           n2181);
   U4599 : AO2 port map( A => n5025, B => n5049, C => n5047, D => n3628, Z => 
                           n3679);
   U4600 : AO2 port map( A => n3665, B => n3340, C => n3328, D => n3666, Z => 
                           n3664);
   U4601 : AO2 port map( A => n3328, B => n3366, C => n2455, D => n3340, Z => 
                           n3398);
   U4602 : AO7 port map( A => n2704, B => n2705, C => n5043, Z => n2703);
   U4603 : AO4 port map( A => n4704, B => n2608, C => n1959, D => n2708, Z => 
                           n2704);
   U4604 : AO4 port map( A => n4705, B => n2706, C => n2707, D => n4687, Z => 
                           n2705);
   U4605 : AO7 port map( A => n4868, B => n2557, C => n4372, Z => n2555);
   U4606 : AO4 port map( A => n4902, B => n4689, C => n4688, D => n2559, Z => 
                           n2557);
   U4607 : AO2 port map( A => n2509, B => n5042, C => n2561, D => n5043, Z => 
                           n2560);
   U4608 : AO7 port map( A => n2538, B => n2539, C => n4371, Z => n2537);
   U4609 : AO4 port map( A => n2541, B => n2542, C => n4893, D => n2544, Z => 
                           n2538);
   U4610 : AO4 port map( A => n4689, B => n2540, C => n4511, D => n4688, Z => 
                           n2539);
   U4611 : AO7 port map( A => n3109, B => n3110, C => n5038, Z => n3108);
   U4612 : AO4 port map( A => n4698, B => n3011, C => n2957, D => n3113, Z => 
                           n3109);
   U4613 : AO4 port map( A => n4700, B => n3111, C => n3112, D => n4682, Z => 
                           n3110);
   U4614 : AO7 port map( A => n4920, B => n2961, C => n4374, Z => n2959);
   U4615 : AO4 port map( A => n4927, B => n4684, C => n4685, D => n2962, Z => 
                           n2961);
   U4616 : AO2 port map( A => n2913, B => n5037, C => n2964, D => n5038, Z => 
                           n2963);
   U4617 : AO7 port map( A => n2944, B => n2945, C => n4369, Z => n2943);
   U4618 : AO4 port map( A => n2946, B => n2947, C => n5068, D => n2949, Z => 
                           n2944);
   U4619 : AO4 port map( A => n4684, B => n1722, C => n4512, D => n4685, Z => 
                           n2945);
   U4620 : AO2 port map( A => n4909, B => n2230, C => n4506, D => n2231, Z => 
                           n2223);
   U4621 : AO3 port map( A => n4972, B => n2236, C => n2237, D => n2238, Z => 
                           n2230);
   U4622 : EO1 port map( A => n4987, B => n4701, C => n2182, D => n4690, Z => 
                           n2233);
   U4623 : AO2 port map( A => n4506, B => n2040, C => n2041, D => n4396, Z => 
                           n2028);
   U4624 : AO4 port map( A => n4359, B => n2047, C => n2048, D => n4361, Z => 
                           n2040);
   U4625 : EON1 port map( A => n4690, B => n2044, C => n4379, D => n2046, Z => 
                           n2041);
   U4626 : AO7 port map( A => n3510, B => n3511, C => n5045, Z => n3509);
   U4627 : AO4 port map( A => n4695, B => n3412, C => n3359, D => n3514, Z => 
                           n3510);
   U4628 : AO4 port map( A => n4697, B => n3512, C => n3513, D => n4678, Z => 
                           n3511);
   U4629 : AO7 port map( A => n5002, B => n3363, C => n4373, Z => n3361);
   U4630 : AO4 port map( A => n5009, B => n4680, C => n4681, D => n3364, Z => 
                           n3363);
   U4631 : AO2 port map( A => n3315, B => n5044, C => n3366, D => n5045, Z => 
                           n3365);
   U4632 : AO7 port map( A => n3346, B => n3347, C => n4370, Z => n3345);
   U4633 : AO4 port map( A => n3348, B => n3349, C => n5073, D => n3351, Z => 
                           n3346);
   U4634 : AO4 port map( A => n4680, B => n2486, C => n4513, D => n4681, Z => 
                           n3347);
   U4635 : AO4 port map( A => n2742, B => n4704, C => n4705, D => n2657, Z => 
                           n2806);
   U4636 : AO4 port map( A => n3146, B => n4698, C => n4700, D => n3062, Z => 
                           n3225);
   U4637 : AO2 port map( A => n4967, B => n4701, C => n4360, D => n2144, Z => 
                           n2257);
   U4638 : EO1 port map( A => n2234, B => n4379, C => n1913, D => n4359, Z => 
                           n2232);
   U4639 : AO4 port map( A => n3547, B => n4695, C => n4697, D => n3464, Z => 
                           n3626);
   U4640 : AO7 port map( A => n4669, B => n4352, C => n1788, Z => n1798);
   U4641 : AO7 port map( A => n4671, B => n4352, C => n1788, Z => n1787);
   U4642 : AO7 port map( A => n4664, B => n4352, C => n1815, Z => n1826);
   U4643 : AO7 port map( A => n4665, B => n4352, C => n1815, Z => n1819);
   U4644 : AO7 port map( A => v_KEY_COLUMN_8_port, B => n4352, C => n1846, Z =>
                           n1889);
   U4645 : AO7 port map( A => n4658, B => n4352, C => n1846, Z => n1863);
   U4646 : AO2 port map( A => n4702, B => n2190, C => n4379, D => n4958, Z => 
                           n2213);
   U4647 : AO2 port map( A => n2215, B => n4701, C => n4983, D => n4360, Z => 
                           n2214);
   U4648 : NR4 port map( A => n1505, B => n1506, C => n1507, D => n1508, Z => 
                           n1504);
   U4649 : ND4 port map( A => n1509, B => n1510, C => n1511, D => n4515, Z => 
                           n1505);
   U4650 : ND3 port map( A => n2590, B => n4362, C => n4686, Z => n2589);
   U4651 : ND3 port map( A => n2454, B => n4363, C => n4679, Z => n3393);
   U4652 : IVDA port map( A => n1949, Y => n4399, Z => n4689);
   U4653 : IVDA port map( A => n2904, Y => n4402, Z => n4684);
   U4654 : IVDA port map( A => n3306, Y => n4400, Z => n4680);
   U4655 : AO6 port map( A => n3070, B => n3081, C => n4698, Z => n3080);
   U4656 : AO6 port map( A => n3472, B => n3483, C => n4695, Z => n3482);
   U4657 : AO4 port map( A => n2590, B => n4704, C => n1959, D => n2738, Z => 
                           n2804);
   U4658 : AO4 port map( A => n1688, B => n4698, C => n2957, D => n3142, Z => 
                           n3223);
   U4659 : AO4 port map( A => n1912, B => n1913, C => n4691, D => n1914, Z => 
                           n1911);
   U4660 : AO4 port map( A => n2454, B => n4695, C => n3359, D => n3543, Z => 
                           n3624);
   U4661 : EO1 port map( A => n5060, B => n2552, C => n2822, D => n2530, Z => 
                           n2855);
   U4662 : EO1 port map( A => n5057, B => n2955, C => n3208, D => n2936, Z => 
                           n3259);
   U4663 : AO7 port map( A => n4378, B => n2153, C => n4506, Z => n2180);
   U4664 : EO1 port map( A => n5051, B => n3357, C => n3609, D => n3338, Z => 
                           n3661);
   U4665 : AO3 port map( A => n4705, B => n2649, C => n4399, D => n2740, Z => 
                           n2722);
   U4666 : AO6 port map( A => n4872, B => n4357, C => n2741, Z => n2740);
   U4667 : AO4 port map( A => n1959, B => n2583, C => n2742, D => n4704, Z => 
                           n2741);
   U4668 : AO6 port map( A => n2565, B => n4399, C => n2567, Z => n2553);
   U4669 : AO4 port map( A => n4688, B => n2568, C => n4881, D => n2541, Z => 
                           n2567);
   U4670 : AO3 port map( A => n4700, B => n3053, C => n4402, D => n3144, Z => 
                           n3126);
   U4671 : AO6 port map( A => n4944, B => n4355, C => n3145, Z => n3144);
   U4672 : AO4 port map( A => n2957, B => n2986, C => n3146, D => n4698, Z => 
                           n3145);
   U4673 : AO6 port map( A => n2968, B => n4402, C => n2969, Z => n2956);
   U4674 : AO4 port map( A => n4685, B => n2970, C => n4942, D => n2946, Z => 
                           n2969);
   U4675 : AO3 port map( A => n4697, B => n3455, C => n4400, D => n3545, Z => 
                           n3527);
   U4676 : AO6 port map( A => n5026, B => n4356, C => n3546, Z => n3545);
   U4677 : AO4 port map( A => n3359, B => n3387, C => n3547, D => n4695, Z => 
                           n3546);
   U4678 : AO6 port map( A => n3370, B => n4400, C => n3371, Z => n3358);
   U4679 : AO4 port map( A => n4681, B => n3372, C => n5024, D => n3348, Z => 
                           n3371);
   U4680 : AO2 port map( A => n2453, B => n2454, C => n2455, D => n4696, Z => 
                           n2452);
   U4681 : AO2 port map( A => n1951, B => n2590, C => n1958, D => n4703, Z => 
                           n2812);
   U4682 : AO2 port map( A => n1687, B => n1688, C => n1689, D => n4699, Z => 
                           n1686);
   U4683 : EON1 port map( A => n2655, B => n4687, C => n2808, D => n4703, Z => 
                           n2807);
   U4684 : EON1 port map( A => n3060, B => n4682, C => n3227, D => n4699, Z => 
                           n3226);
   U4685 : EON1 port map( A => n3462, B => n4678, C => n3628, D => n4696, Z => 
                           n3627);
   U4686 : AO3 port map( A => n4921, B => n2957, C => n4402, D => n3077, Z => 
                           n3075);
   U4687 : AO3 port map( A => n5003, B => n3359, C => n4400, D => n3479, Z => 
                           n3477);
   U4688 : AO6 port map( A => n2665, B => n2676, C => n4704, Z => n2675);
   U4689 : AO2 port map( A => n4955, B => n4378, C => n4995, D => n4701, Z => 
                           n2253);
   U4690 : AO4 port map( A => n4704, B => n2728, C => n1959, D => n1988, Z => 
                           n2727);
   U4691 : AO4 port map( A => n4698, B => n3132, C => n2957, D => n1713, Z => 
                           n3131);
   U4692 : AO4 port map( A => n4695, B => n3533, C => n3359, D => n2477, Z => 
                           n3532);
   U4693 : AO3 port map( A => n4886, B => n1959, C => n4399, D => n2672, Z => 
                           n2670);
   U4694 : ND3 port map( A => n4873, B => n4368, C => n5043, Z => n2554);
   U4695 : ND3 port map( A => n4950, B => n4364, C => n5038, Z => n2958);
   U4696 : ND3 port map( A => n5032, B => n4367, C => n5045, Z => n3360);
   U4697 : NR3 port map( A => n1498, B => v_CALCULATION_CNTR_3_port, C => n2866
                           , Z => n1351);
   U4698 : NR3 port map( A => v_CALCULATION_CNTR_0_port, B => 
                           v_CALCULATION_CNTR_3_port, C => n1498, Z => n3671);
   U4699 : AO4 port map( A => n4712, B => n297, C => n4383, D => n298, Z => 
                           n296);
   U4700 : AO4 port map( A => n4712, B => n1108, C => n4383, D => n1109, Z => 
                           n1107);
   U4701 : AO3 port map( A => n4354, B => n4464, C => n1319, D => n1320, Z => 
                           n3971);
   U4702 : AO2 port map( A => n1364, B => n1365, C => n4741, D => n1366, Z => 
                           n1319);
   U4703 : AO3 port map( A => n4354, B => n4465, C => n966, D => n967, Z => 
                           n3977);
   U4704 : AO2 port map( A => n4733, B => n994, C => n995, D => n996, Z => n966
                           );
   U4705 : AO3 port map( A => n4354, B => n4466, C => n145, D => n146, Z => 
                           n3983);
   U4706 : AO2 port map( A => n4794, B => n188, C => n189, D => n190, Z => n145
                           );
   U4707 : IVDA port map( A => v_KEY_COLUMN_13_port, Y => n4385, Z => n4660);
   U4708 : IVDA port map( A => v_KEY_COLUMN_5_port, Y => n4461, Z => n4655);
   U4709 : AO4 port map( A => n4712, B => n600, C => n4383, D => n601, Z => 
                           n599);
   U4710 : AO4 port map( A => n4712, B => n429, C => n4383, D => n430, Z => 
                           n428);
   U4711 : AO4 port map( A => n4712, B => n470, C => n4383, D => n471, Z => 
                           n469);
   U4712 : AO4 port map( A => n4712, B => n1069, C => n4383, D => n1070, Z => 
                           n1068);
   U4713 : AO4 port map( A => n4712, B => n735, C => n4383, D => n736, Z => 
                           n734);
   U4714 : AO4 port map( A => n4712, B => n239, C => n4383, D => n240, Z => 
                           n238);
   U4715 : AO4 port map( A => n4712, B => n210, C => n4383, D => n211, Z => 
                           n209);
   U4716 : AO4 port map( A => n4712, B => n1011, C => n4383, D => n1012, Z => 
                           n1010);
   U4717 : AO4 port map( A => v_RAM_OUT0_9_port, B => n1890, C => n2393, D => 
                           n4569, Z => n1558);
   U4718 : AO4 port map( A => n4690, B => n1913, C => n4956, D => n4361, Z => 
                           n2394);
   U4719 : AO6 port map( A => n2396, B => n2397, C => v_RAM_OUT0_15_port, Z => 
                           n2395);
   U4720 : ND3 port map( A => n1350, B => n4354, C => n1351, Z => n164);
   U4721 : IVDA port map( A => v_KEY_COLUMN_22_port, Y => n4460, Z => n4665);
   U4722 : IVDA port map( A => v_KEY_COLUMN_23_port, Y => n4387, Z => n4666);
   U4723 : IVDA port map( A => v_KEY_COLUMN_15_port, Y => n4388, Z => n4662);
   U4724 : AO3 port map( A => n1558, B => n2020, C => n2388, D => n2389, Z => 
                           n4174);
   U4725 : AO7 port map( A => v_KEY_COLUMN_8_port, B => n4706, C => n2024, Z =>
                           n2390);
   U4726 : AO3 port map( A => n1523, B => n1558, C => n1559, D => n1560, Z => 
                           n4206);
   U4727 : AO7 port map( A => v_KEY_COLUMN_8_port, B => n1527, C => n1529, Z =>
                           n1561);
   U4728 : AO3 port map( A => n1558, B => n1726, C => n1751, D => n1752, Z => 
                           n4238);
   U4729 : AO7 port map( A => v_KEY_COLUMN_8_port, B => n1609, C => n1731, Z =>
                           n1753);
   U4730 : IVDA port map( A => v_KEY_COLUMN_30_port, Y => n4573, Z => n4670);
   U4731 : IVDA port map( A => v_KEY_COLUMN_31_port, Y => n4459, Z => n4671);
   U4732 : IVDA port map( A => v_KEY_COLUMN_14_port, Y => n4577, Z => n4661);
   U4733 : IVDA port map( A => v_KEY_COLUMN_6_port, Y => n4574, Z => n4656);
   U4734 : IVDA port map( A => v_KEY_COLUMN_7_port, Y => n4575, Z => n4657);
   U4735 : IVDA port map( A => v_KEY_COLUMN_10_port, Y => n4390, Z => n4658);
   U4736 : AO3 port map( A => n1886, B => n1841, C => n1887, D => n1888, Z => 
                           n4270);
   U4737 : AO6 port map( A => n1890, B => n4569, C => n1892, Z => n1886);
   U4738 : AO4 port map( A => n2975, B => n2976, C => n2977, D => n4578, Z => 
                           n1651);
   U4739 : AO3 port map( A => n3030, B => n2949, C => n3031, D => n4578, Z => 
                           n2975);
   U4740 : AO2 port map( A => v_RAM_OUT0_21_port, B => n2978, C => n2979, D => 
                           n4409, Z => n2977);
   U4741 : AO7 port map( A => n4852, B => n4463, C => n1477, Z => n1475);
   U4742 : IVDA port map( A => v_KEY_COLUMN_24_port, Y => n4571, Z => n4667);
   U4743 : IVDA port map( A => v_KEY_COLUMN_27_port, Y => n4572, Z => n4668);
   U4744 : IVDA port map( A => v_KEY_COLUMN_28_port, Y => n4458, Z => n4669);
   U4745 : IVDA port map( A => v_KEY_COLUMN_17_port, Y => n4403, Z => n4663);
   U4746 : AO2 port map( A => n5039, B => n1902, C => v_RAM_OUT0_13_port, D => 
                           n2398, Z => n2397);
   U4747 : AO7 port map( A => n5064, B => n4975, C => n2401, Z => n2398);
   U4748 : AO2 port map( A => n4701, B => n4974, C => n4980, D => n4360, Z => 
                           n2401);
   U4749 : AO3 port map( A => n1640, B => n1917, C => n1963, D => n1964, Z => 
                           n4032);
   U4750 : AO7 port map( A => n4667, B => n4706, C => n1923, Z => n1965);
   U4751 : AO3 port map( A => n1636, B => n1917, C => n1960, D => n1961, Z => 
                           n4075);
   U4752 : AO7 port map( A => v_KEY_COLUMN_25_port, B => n4706, C => n1923, Z 
                           => n1962);
   U4753 : AO3 port map( A => n1632, B => n1917, C => n1938, D => n1939, Z => 
                           n4106);
   U4754 : AO7 port map( A => v_KEY_COLUMN_26_port, B => n4706, C => n1923, Z 
                           => n1940);
   U4755 : AO3 port map( A => n1627, B => n1917, C => n1935, D => n1936, Z => 
                           n4131);
   U4756 : AO7 port map( A => n4668, B => n4706, C => n1923, Z => n1937);
   U4757 : AO3 port map( A => n1612, B => n1917, C => n1924, D => n1925, Z => 
                           n4164);
   U4758 : AO7 port map( A => n4670, B => n4706, C => n1923, Z => n1926);
   U4759 : AO3 port map( A => n1837, B => n1991, C => n2015, D => n2016, Z => 
                           n4166);
   U4760 : AO7 port map( A => v_KEY_COLUMN_16_port, B => n4706, C => n1995, Z 
                           => n2017);
   U4761 : AO3 port map( A => n1694, B => n1991, C => n2012, D => n2013, Z => 
                           n4167);
   U4762 : AO7 port map( A => n4663, B => n4706, C => n1995, Z => n2014);
   U4763 : AO3 port map( A => n1830, B => n1991, C => n2009, D => n2010, Z => 
                           n4168);
   U4764 : AO7 port map( A => v_KEY_COLUMN_18_port, B => n4706, C => n1995, Z 
                           => n2011);
   U4765 : AO3 port map( A => n1667, B => n1991, C => n2006, D => n2007, Z => 
                           n4169);
   U4766 : AO7 port map( A => v_KEY_COLUMN_19_port, B => n4706, C => n1995, Z 
                           => n2008);
   U4767 : AO3 port map( A => n1661, B => n1991, C => n2002, D => n2003, Z => 
                           n4170);
   U4768 : AO7 port map( A => n4664, B => n4706, C => n1995, Z => n2005);
   U4769 : AO3 port map( A => n1645, B => n1991, C => n1992, D => n1993, Z => 
                           n4173);
   U4770 : AO7 port map( A => n4666, B => n4706, C => n1995, Z => n1994);
   U4771 : EON1 port map( A => n4619, B => n1476, C => n4619, D => n1475, Z => 
                           n4287);
   U4772 : AO4 port map( A => n2573, B => n2574, C => n2575, D => n4587, Z => 
                           n1612);
   U4773 : AO3 port map( A => n2626, B => n2544, C => n2627, D => n4587, Z => 
                           n2573);
   U4774 : AO2 port map( A => v_RAM_OUT0_29_port, B => n2576, C => n2577, D => 
                           n4410, Z => n2575);
   U4775 : AO4 port map( A => n2496, B => n2497, C => v_RAM_OUT0_31_port, D => 
                           n2498, Z => n1603);
   U4776 : AO3 port map( A => n2536, B => n4687, C => n2537, D => 
                           v_RAM_OUT0_31_port, Z => n2497);
   U4777 : AO3 port map( A => n2553, B => n1959, C => n2554, D => n2555, Z => 
                           n2496);
   U4778 : AO6 port map( A => v_RAM_OUT0_29_port, B => n2499, C => n2500, Z => 
                           n2498);
   U4779 : AO4 port map( A => n2898, B => n2899, C => v_RAM_OUT0_23_port, D => 
                           n2900, Z => n1645);
   U4780 : AO3 port map( A => n2942, B => n4682, C => n2943, D => 
                           v_RAM_OUT0_23_port, Z => n2899);
   U4781 : AO3 port map( A => n2956, B => n2957, C => n2958, D => n2959, Z => 
                           n2898);
   U4782 : AO6 port map( A => v_RAM_OUT0_21_port, B => n2901, C => n2902, Z => 
                           n2900);
   U4783 : AO4 port map( A => n2353, B => n4569, C => v_RAM_OUT0_9_port, D => 
                           n2354, Z => n1553);
   U4784 : AO6 port map( A => v_RAM_OUT0_15_port, B => n2373, C => n2374, Z => 
                           n2353);
   U4785 : AO6 port map( A => v_RAM_OUT0_15_port, B => n2355, C => n2356, Z => 
                           n2354);
   U4786 : AO4 port map( A => n2375, B => n1897, C => n2376, D => n4691, Z => 
                           n2374);
   U4787 : AO3 port map( A => n2269, B => n4569, C => n2270, D => n2271, Z => 
                           n1544);
   U4788 : ND4 port map( A => n2272, B => n4904, C => n2274, D => n2275, Z => 
                           n2271);
   U4789 : ND4 port map( A => n2285, B => n4907, C => n2286, D => n2287, Z => 
                           n2270);
   U4790 : AO6 port map( A => v_RAM_OUT0_15_port, B => n2296, C => n2297, Z => 
                           n2269);
   U4791 : AO4 port map( A => v_RAM_OUT0_9_port, B => n2171, C => n2172, D => 
                           n4569, Z => n1535);
   U4792 : AO7 port map( A => v_RAM_OUT0_9_port, B => n2025, C => n2026, Z => 
                           n1522);
   U4793 : ND4 port map( A => v_RAM_OUT0_9_port, B => n2027, C => n2028, D => 
                           n2029, Z => n2026);
   U4794 : AO4 port map( A => n3376, B => n3377, C => n3378, D => n4588, Z => 
                           n1570);
   U4795 : AO3 port map( A => n3431, B => n3351, C => n3432, D => n4588, Z => 
                           n3376);
   U4796 : AO2 port map( A => v_RAM_OUT0_5_port, B => n3379, C => n3380, D => 
                           n4408, Z => n3378);
   U4797 : AO4 port map( A => n3300, B => n3301, C => v_RAM_OUT0_7_port, D => 
                           n3302, Z => n1563);
   U4798 : AO3 port map( A => n3344, B => n4678, C => n3345, D => 
                           v_RAM_OUT0_7_port, Z => n3301);
   U4799 : AO3 port map( A => n3358, B => n3359, C => n3360, D => n3361, Z => 
                           n3300);
   U4800 : AO6 port map( A => v_RAM_OUT0_5_port, B => n3303, C => n3304, Z => 
                           n3302);
   U4801 : AO4 port map( A => n1966, B => n4587, C => v_RAM_OUT0_31_port, D => 
                           n1967, Z => n1640);
   U4802 : AO2 port map( A => n1968, B => n1969, C => n1970, D => n4410, Z => 
                           n1967);
   U4803 : AO6 port map( A => v_RAM_OUT0_29_port, B => n1982, C => n1983, Z => 
                           n1966);
   U4804 : AO6 port map( A => n1980, B => n4499, C => n4410, Z => n1968);
   U4805 : AO4 port map( A => n3269, B => n4578, C => v_RAM_OUT0_23_port, D => 
                           n3270, Z => n1837);
   U4806 : AO2 port map( A => n3271, B => n3272, C => n1716, D => n4409, Z => 
                           n3270);
   U4807 : AO6 port map( A => v_RAM_OUT0_21_port, B => n1705, C => n3281, Z => 
                           n3269);
   U4808 : AO6 port map( A => n1720, B => n4498, C => n4409, Z => n3271);
   U4809 : AO4 port map( A => n3673, B => n4588, C => v_RAM_OUT0_7_port, D => 
                           n3674, Z => n1598);
   U4810 : AO2 port map( A => n3675, B => n3676, C => n2480, D => n4408, Z => 
                           n3674);
   U4811 : AO6 port map( A => v_RAM_OUT0_5_port, B => n2469, C => n3685, Z => 
                           n3673);
   U4812 : AO6 port map( A => n2484, B => n4497, C => n4408, Z => n3675);
   U4813 : ND4 port map( A => v_RAM_OUT0_9_port, B => n2222, C => n2223, D => 
                           n2224, Z => n2221);
   U4814 : AO3 port map( A => n2247, B => n1912, C => n2248, D => n2249, Z => 
                           n2220);
   U4815 : IVDA port map( A => n1724, Y => n4512, Z => n4683);
   U4816 : IVDA port map( A => n2488, Y => n4513, Z => n4679);
   U4817 : IVDA port map( A => n1483, Y => n4565, Z => n4672);
   U4818 : AO3 port map( A => n2318, B => n2178, C => n2319, D => n2320, Z => 
                           n1869);
   U4819 : AO2 port map( A => n5040, B => n2325, C => n2032, D => n2054, Z => 
                           n2319);
   U4820 : AO2 port map( A => v_RAM_OUT0_13_port, B => n2321, C => n2065, D => 
                           n2290, Z => n2320);
   U4821 : AO6 port map( A => n2252, B => n2253, C => n2074, Z => n2251);
   U4822 : AO2 port map( A => n2145, B => n4702, C => n4966, D => n4379, Z => 
                           n2256);
   U4823 : IVDA port map( A => v_KEY_COLUMN_20_port, Y => n4457, Z => n4664);
   U4824 : IVDA port map( A => v_KEY_COLUMN_11_port, Y => n4576, Z => n4659);
   U4825 : AO4 port map( A => n3044, B => n3045, C => v_RAM_OUT0_23_port, D => 
                           n3046, Z => n3043);
   U4826 : AO4 port map( A => n3446, B => n3447, C => v_RAM_OUT0_7_port, D => 
                           n3448, Z => n3445);
   U4827 : EON1 port map( A => n2529, B => n2530, C => n4889, D => n2531, Z => 
                           n2516);
   U4828 : AO4 port map( A => n2533, B => n2534, C => v_RAM_OUT0_25_port, D => 
                           n4879, Z => n2515);
   U4829 : AO3 port map( A => n4872, B => n2519, C => n2520, D => n2521, Z => 
                           n2517);
   U4830 : EON1 port map( A => n2935, B => n2936, C => n4949, D => n2938, Z => 
                           n2920);
   U4831 : AO4 port map( A => n2939, B => n2940, C => v_RAM_OUT0_17_port, D => 
                           n4923, Z => n2919);
   U4832 : AO3 port map( A => n4944, B => n2923, C => n2924, D => n2925, Z => 
                           n2921);
   U4833 : EON1 port map( A => n3337, B => n3338, C => n5031, D => n3340, Z => 
                           n3322);
   U4834 : AO4 port map( A => n3341, B => n3342, C => v_RAM_OUT0_1_port, D => 
                           n5005, Z => n3321);
   U4835 : AO3 port map( A => n5026, B => n3325, C => n3326, D => n3327, Z => 
                           n3323);
   U4836 : AO2 port map( A => n3072, B => n4683, C => n4941, D => 
                           v_RAM_OUT0_20_port, Z => n3071);
   U4837 : AO2 port map( A => n3474, B => n4679, C => n5023, D => 
                           v_RAM_OUT0_4_port, Z => n3473);
   U4838 : EO1 port map( A => v_RAM_OUT0_25_port, B => n2882, C => n2619, D => 
                           n2519, Z => n2881);
   U4839 : AO3 port map( A => n4362, B => n2586, C => n4879, D => n2883, Z => 
                           n2882);
   U4840 : EO1 port map( A => n4878, B => v_RAM_OUT0_28_port, C => n1959, D => 
                           n2655, Z => n2883);
   U4841 : EO1 port map( A => v_RAM_OUT0_17_port, B => n3293, C => n3022, D => 
                           n2923, Z => n3292);
   U4842 : AO3 port map( A => n4365, B => n2989, C => n4923, D => n3294, Z => 
                           n3293);
   U4843 : EO1 port map( A => n4940, B => v_RAM_OUT0_20_port, C => n2957, D => 
                           n3060, Z => n3294);
   U4844 : EO1 port map( A => v_RAM_OUT0_1_port, B => n3697, C => n3423, D => 
                           n3325, Z => n3696);
   U4845 : AO3 port map( A => n4363, B => n3390, C => n5005, D => n3698, Z => 
                           n3697);
   U4846 : EO1 port map( A => n5022, B => v_RAM_OUT0_4_port, C => n3359, D => 
                           n3462, Z => n3698);
   U4847 : AO7 port map( A => n3032, B => n3033, C => n5037, Z => n3031);
   U4848 : AO3 port map( A => n4945, B => n2957, C => n3034, D => n3028, Z => 
                           n3032);
   U4849 : AO4 port map( A => n1725, B => n4698, C => v_RAM_OUT0_20_port, D => 
                           n2965, Z => n3033);
   U4850 : AO3 port map( A => n2363, B => n4516, C => n2364, D => n2365, Z => 
                           n2355);
   U4851 : AO2 port map( A => n5041, B => n2212, C => n2065, D => n4992, Z => 
                           n2365);
   U4852 : AO2 port map( A => n2367, B => v_RAM_OUT0_10_port, C => n2054, D => 
                           n2072, Z => n2364);
   U4853 : AO3 port map( A => n2383, B => n4516, C => n2384, D => n2385, Z => 
                           n2373);
   U4854 : AO2 port map( A => n2386, B => n2065, C => n2054, D => n2192, Z => 
                           n2384);
   U4855 : AO2 port map( A => n5040, B => n2038, C => n5041, D => n1900, Z => 
                           n2385);
   U4856 : AO3 port map( A => n2306, B => n2183, C => n2307, D => n2308, Z => 
                           n2296);
   U4857 : AO2 port map( A => n2065, B => n1900, C => n5041, D => n4971, Z => 
                           n2308);
   U4858 : AO2 port map( A => v_RAM_OUT0_13_port, B => n2309, C => n2054, D => 
                           n4959, Z => n2307);
   U4859 : AO3 port map( A => n4971, B => n2227, C => n2311, D => n2312, Z => 
                           n2309);
   U4860 : AO3 port map( A => n2129, B => n2183, C => n2184, D => n2185, Z => 
                           n2173);
   U4861 : AO2 port map( A => n2065, B => n2186, C => n2159, D => n5041, Z => 
                           n2185);
   U4862 : AO2 port map( A => n2113, B => n2054, C => v_RAM_OUT0_13_port, D => 
                           n2187, Z => n2184);
   U4863 : ND4 port map( A => n2123, B => v_RAM_OUT0_15_port, C => n2124, D => 
                           n2125, Z => n2106);
   U4864 : AO2 port map( A => n2131, B => n2065, C => n4961, D => n2054, Z => 
                           n2124);
   U4865 : AO7 port map( A => n2126, B => n2127, C => v_RAM_OUT0_13_port, Z => 
                           n2125);
   U4866 : AO2 port map( A => n4989, B => n5040, C => n5041, D => n1900, Z => 
                           n2123);
   U4867 : AO4 port map( A => n1866, B => n1867, C => n1868, D => n1869, Z => 
                           n1865);
   U4868 : AO3 port map( A => n1876, B => n1877, C => n1878, D => n1879, Z => 
                           n1866);
   U4869 : AO3 port map( A => n1870, B => n4516, C => n1872, D => n4907, Z => 
                           n1867);
   U4870 : AO7 port map( A => v_RAM_OUT0_31_port, B => n2827, C => n2828, Z => 
                           n1636);
   U4871 : AO6 port map( A => v_RAM_OUT0_29_port, B => n2843, C => n2844, Z => 
                           n2827);
   U4872 : AO3 port map( A => n2829, B => n2830, C => v_RAM_OUT0_31_port, D => 
                           n2831, Z => n2828);
   U4873 : ND4 port map( A => n2855, B => n2856, C => n2857, D => n2858, Z => 
                           n2843);
   U4874 : AO7 port map( A => v_RAM_OUT0_23_port, B => n3231, C => n3232, Z => 
                           n1694);
   U4875 : AO6 port map( A => v_RAM_OUT0_21_port, B => n3247, C => n3248, Z => 
                           n3231);
   U4876 : AO3 port map( A => n3233, B => n3234, C => v_RAM_OUT0_23_port, D => 
                           n3235, Z => n3232);
   U4877 : ND4 port map( A => n3259, B => n3260, C => n3261, D => n3262, Z => 
                           n3247);
   U4878 : AO7 port map( A => v_RAM_OUT0_9_port, B => n2104, C => n2105, Z => 
                           n1530);
   U4879 : ND4 port map( A => v_RAM_OUT0_9_port, B => n2106, C => n2107, D => 
                           n2108, Z => n2105);
   U4880 : AO6 port map( A => v_RAM_OUT0_15_port, B => n2136, C => n2137, Z => 
                           n2104);
   U4881 : AO3 port map( A => n4359, B => n2064, C => n4906, D => n2117, Z => 
                           n2107);
   U4882 : AO7 port map( A => v_RAM_OUT0_7_port, B => n3633, C => n3634, Z => 
                           n1593);
   U4883 : AO6 port map( A => v_RAM_OUT0_5_port, B => n3649, C => n3650, Z => 
                           n3633);
   U4884 : AO3 port map( A => n3635, B => n3636, C => v_RAM_OUT0_7_port, D => 
                           n3637, Z => n3634);
   U4885 : ND4 port map( A => n3661, B => n3662, C => n3663, D => n3664, Z => 
                           n3649);
   U4886 : AO6 port map( A => n3063, B => n3064, C => n4409, Z => n3047);
   U4887 : AO2 port map( A => v_RAM_OUT0_17_port, B => n3068, C => n4948, D => 
                           n5055, Z => n3063);
   U4888 : AO3 port map( A => n1725, B => n4700, C => n3065, D => n3066, Z => 
                           n3064);
   U4889 : AO4 port map( A => n4365, B => n3070, C => v_RAM_OUT0_18_port, D => 
                           n3071, Z => n3068);
   U4890 : AO6 port map( A => n3465, B => n3466, C => n4408, Z => n3449);
   U4891 : AO2 port map( A => v_RAM_OUT0_1_port, B => n3470, C => n5030, D => 
                           n5049, Z => n3465);
   U4892 : AO3 port map( A => n2489, B => n4697, C => n3467, D => n3468, Z => 
                           n3466);
   U4893 : AO4 port map( A => n4363, B => n3472, C => v_RAM_OUT0_2_port, D => 
                           n3473, Z => n3470);
   U4894 : AO3 port map( A => n1553, B => n2020, C => n2350, D => n2351, Z => 
                           n4175);
   U4895 : AO7 port map( A => v_KEY_COLUMN_9_port, B => n4706, C => n2024, Z =>
                           n2352);
   U4896 : AO3 port map( A => n1549, B => n2020, C => n2313, D => n2314, Z => 
                           n4176);
   U4897 : AO7 port map( A => n4658, B => n4706, C => n2024, Z => n2315);
   U4898 : AO3 port map( A => n1544, B => n2020, C => n2266, D => n2267, Z => 
                           n4177);
   U4899 : AO7 port map( A => n4659, B => n4706, C => n2024, Z => n2268);
   U4900 : AO3 port map( A => n1540, B => n2020, C => n2217, D => n2218, Z => 
                           n4178);
   U4901 : AO7 port map( A => v_KEY_COLUMN_12_port, B => n4706, C => n2024, Z 
                           => n2219);
   U4902 : AO3 port map( A => n1535, B => n2020, C => n2168, D => n2169, Z => 
                           n4179);
   U4903 : AO7 port map( A => n4660, B => n4706, C => n2024, Z => n2170);
   U4904 : AO3 port map( A => n1530, B => n2020, C => n2101, D => n2102, Z => 
                           n4180);
   U4905 : AO7 port map( A => n4661, B => n4706, C => n2024, Z => n2103);
   U4906 : AO3 port map( A => n1522, B => n2020, C => n2021, D => n2022, Z => 
                           n4181);
   U4907 : AO7 port map( A => n4662, B => n4706, C => n2024, Z => n2023);
   U4908 : AO3 port map( A => n2463, B => n2422, C => n2464, D => n2465, Z => 
                           n4182);
   U4909 : AO2 port map( A => n2467, B => n4588, C => v_RAM_OUT0_7_port, D => 
                           n2468, Z => n2463);
   U4910 : AO3 port map( A => n1593, B => n2422, C => n2460, D => n2461, Z => 
                           n4183);
   U4911 : AO7 port map( A => v_KEY_COLUMN_1_port, B => n4706, C => n2426, Z =>
                           n2462);
   U4912 : AO3 port map( A => n2437, B => n2422, C => n2438, D => n2439, Z => 
                           n4184);
   U4913 : AO2 port map( A => v_RAM_OUT0_7_port, B => n2441, C => n5004, D => 
                           n4588, Z => n2437);
   U4914 : AO3 port map( A => n1585, B => n2422, C => n2434, D => n2435, Z => 
                           n4185);
   U4915 : AO7 port map( A => v_KEY_COLUMN_3_port, B => n4706, C => n2426, Z =>
                           n2436);
   U4916 : AO3 port map( A => n1581, B => n2422, C => n2431, D => n2432, Z => 
                           n4186);
   U4917 : AO7 port map( A => v_KEY_COLUMN_4_port, B => n4706, C => n2426, Z =>
                           n2433);
   U4918 : AO3 port map( A => n1570, B => n2422, C => n2427, D => n2428, Z => 
                           n4188);
   U4919 : AO7 port map( A => n4656, B => n4706, C => n2426, Z => n2429);
   U4920 : AO3 port map( A => n1563, B => n2422, C => n2423, D => n2424, Z => 
                           n4189);
   U4921 : AO7 port map( A => n4657, B => n4706, C => n2426, Z => n2425);
   U4922 : AO3 port map( A => n2862, B => n2490, C => n2863, D => n2864, Z => 
                           n4190);
   U4923 : AO2 port map( A => n2867, B => n4587, C => v_RAM_OUT0_31_port, D => 
                           n2868, Z => n2862);
   U4924 : AO3 port map( A => n1636, B => n2490, C => n2824, D => n2825, Z => 
                           n4191);
   U4925 : AO7 port map( A => v_KEY_COLUMN_25_port, B => n1527, C => n2495, Z 
                           => n2826);
   U4926 : AO3 port map( A => n2787, B => n2490, C => n2788, D => n2789, Z => 
                           n4192);
   U4927 : AO2 port map( A => v_RAM_OUT0_31_port, B => n2791, C => n4867, D => 
                           n4587, Z => n2787);
   U4928 : AO3 port map( A => n1627, B => n2490, C => n2743, D => n2744, Z => 
                           n4193);
   U4929 : AO7 port map( A => n4668, B => n1527, C => n2495, Z => n2745);
   U4930 : AO3 port map( A => n1621, B => n2490, C => n2695, D => n2696, Z => 
                           n4194);
   U4931 : AO7 port map( A => n4669, B => n1527, C => n2495, Z => n2698);
   U4932 : AO3 port map( A => n4870, B => n2490, C => n2636, D => n2637, Z => 
                           n4195);
   U4933 : AO7 port map( A => v_KEY_COLUMN_29_port, B => n1527, C => n2495, Z 
                           => n2638);
   U4934 : AO3 port map( A => n1612, B => n2490, C => n2570, D => n2571, Z => 
                           n4196);
   U4935 : AO7 port map( A => n4670, B => n1527, C => n2495, Z => n2572);
   U4936 : AO3 port map( A => n1603, B => n2490, C => n2491, D => n2492, Z => 
                           n4197);
   U4937 : AO7 port map( A => n4671, B => n1527, C => n2495, Z => n2494);
   U4938 : AO3 port map( A => n1837, B => n2893, C => n3266, D => n3267, Z => 
                           n4198);
   U4939 : AO7 port map( A => v_KEY_COLUMN_16_port, B => n1527, C => n2897, Z 
                           => n3268);
   U4940 : AO3 port map( A => n1694, B => n2893, C => n3228, D => n3229, Z => 
                           n4199);
   U4941 : AO7 port map( A => n4663, B => n1527, C => n2897, Z => n3230);
   U4942 : AO3 port map( A => n1830, B => n2893, C => n3192, D => n3193, Z => 
                           n4200);
   U4943 : AO7 port map( A => v_KEY_COLUMN_18_port, B => n1527, C => n2897, Z 
                           => n3194);
   U4944 : AO3 port map( A => n1667, B => n2893, C => n3147, D => n3148, Z => 
                           n4201);
   U4945 : AO7 port map( A => v_KEY_COLUMN_19_port, B => n1527, C => n2897, Z 
                           => n3149);
   U4946 : AO3 port map( A => n4903, B => n2893, C => n3040, D => n3041, Z => 
                           n4203);
   U4947 : AO7 port map( A => v_KEY_COLUMN_21_port, B => n1527, C => n2897, Z 
                           => n3042);
   U4948 : AO3 port map( A => n1645, B => n2893, C => n2894, D => n2895, Z => 
                           n4205);
   U4949 : AO7 port map( A => n4666, B => n1527, C => n2897, Z => n2896);
   U4950 : AO3 port map( A => n1523, B => n1553, C => n1554, D => n1555, Z => 
                           n4207);
   U4951 : AO7 port map( A => v_KEY_COLUMN_9_port, B => n1527, C => n1529, Z =>
                           n1557);
   U4952 : AO3 port map( A => n1523, B => n1549, C => n1550, D => n1551, Z => 
                           n4208);
   U4953 : AO7 port map( A => n4658, B => n1527, C => n1529, Z => n1552);
   U4954 : AO3 port map( A => n1523, B => n1544, C => n1545, D => n1546, Z => 
                           n4209);
   U4955 : AO7 port map( A => n4659, B => n1527, C => n1529, Z => n1548);
   U4956 : AO3 port map( A => n1523, B => n1540, C => n1541, D => n1542, Z => 
                           n4210);
   U4957 : AO7 port map( A => v_KEY_COLUMN_12_port, B => n1527, C => n1529, Z 
                           => n1543);
   U4958 : AO3 port map( A => n1523, B => n1535, C => n1536, D => n1537, Z => 
                           n4211);
   U4959 : AO7 port map( A => n4660, B => n1527, C => n1529, Z => n1539);
   U4960 : AO3 port map( A => n1523, B => n1530, C => n1531, D => n1532, Z => 
                           n4212);
   U4961 : AO7 port map( A => n4661, B => n1527, C => n1529, Z => n1534);
   U4962 : AO3 port map( A => n1522, B => n1523, C => n1524, D => n1525, Z => 
                           n4213);
   U4963 : AO7 port map( A => n4662, B => n1527, C => n1529, Z => n1528);
   U4964 : AO3 port map( A => n1564, B => n1598, C => n1599, D => n1600, Z => 
                           n4214);
   U4965 : AO7 port map( A => v_KEY_COLUMN_0_port, B => n1527, C => n1569, Z =>
                           n1601);
   U4966 : AO3 port map( A => n1564, B => n1593, C => n1594, D => n1595, Z => 
                           n4215);
   U4967 : AO7 port map( A => v_KEY_COLUMN_1_port, B => n1527, C => n1569, Z =>
                           n1597);
   U4968 : AO3 port map( A => n1564, B => n1589, C => n1590, D => n1591, Z => 
                           n4216);
   U4969 : AO7 port map( A => v_KEY_COLUMN_2_port, B => n1527, C => n1569, Z =>
                           n1592);
   U4970 : AO3 port map( A => n1564, B => n1585, C => n1586, D => n1587, Z => 
                           n4217);
   U4971 : AO7 port map( A => v_KEY_COLUMN_3_port, B => n1527, C => n1569, Z =>
                           n1588);
   U4972 : AO3 port map( A => n1564, B => n1581, C => n1582, D => n1583, Z => 
                           n4218);
   U4973 : AO7 port map( A => v_KEY_COLUMN_4_port, B => n1527, C => n1569, Z =>
                           n1584);
   U4974 : AO3 port map( A => n4911, B => n1564, C => n1576, D => n1577, Z => 
                           n4219);
   U4975 : AO7 port map( A => n4655, B => n1527, C => n1569, Z => n1580);
   U4976 : AO3 port map( A => n1564, B => n1570, C => n1571, D => n1572, Z => 
                           n4220);
   U4977 : AO7 port map( A => n4656, B => n1527, C => n1569, Z => n1574);
   U4978 : AO3 port map( A => n1563, B => n1564, C => n1565, D => n1566, Z => 
                           n4221);
   U4979 : AO7 port map( A => n4657, B => n1527, C => n1569, Z => n1568);
   U4980 : AO3 port map( A => n1604, B => n1640, C => n1641, D => n1642, Z => 
                           n4222);
   U4981 : AO7 port map( A => n4667, B => n1609, C => n1611, Z => n1644);
   U4982 : AO3 port map( A => n1604, B => n1636, C => n1637, D => n1638, Z => 
                           n4223);
   U4983 : AO7 port map( A => v_KEY_COLUMN_25_port, B => n1609, C => n1611, Z 
                           => n1639);
   U4984 : AO3 port map( A => n1604, B => n1632, C => n1633, D => n1634, Z => 
                           n4224);
   U4985 : AO7 port map( A => v_KEY_COLUMN_26_port, B => n1609, C => n1611, Z 
                           => n1635);
   U4986 : AO3 port map( A => n1604, B => n1627, C => n1628, D => n1629, Z => 
                           n4225);
   U4987 : AO7 port map( A => n4668, B => n1609, C => n1611, Z => n1631);
   U4988 : AO3 port map( A => n1604, B => n1621, C => n1622, D => n1623, Z => 
                           n4226);
   U4989 : AO7 port map( A => n4669, B => n1609, C => n1611, Z => n1626);
   U4990 : AO3 port map( A => n4870, B => n1604, C => n1618, D => n1619, Z => 
                           n4227);
   U4991 : AO7 port map( A => v_KEY_COLUMN_29_port, B => n1609, C => n1611, Z 
                           => n1620);
   U4992 : AO3 port map( A => n1604, B => n1612, C => n1613, D => n1614, Z => 
                           n4228);
   U4993 : AO7 port map( A => n4670, B => n1609, C => n1611, Z => n1616);
   U4994 : AO3 port map( A => n1603, B => n1604, C => n1605, D => n1606, Z => 
                           n4229);
   U4995 : AO7 port map( A => n4671, B => n1609, C => n1611, Z => n1610);
   U4996 : AO3 port map( A => n1698, B => n1646, C => n1699, D => n1700, Z => 
                           n4230);
   U4997 : AO2 port map( A => n1703, B => n4578, C => v_RAM_OUT0_23_port, D => 
                           n1704, Z => n1698);
   U4998 : AO3 port map( A => n1646, B => n1694, C => n1695, D => n1696, Z => 
                           n4231);
   U4999 : AO7 port map( A => n4663, B => n1609, C => n1650, Z => n1697);
   U5000 : AO3 port map( A => n1671, B => n1646, C => n1672, D => n1673, Z => 
                           n4232);
   U5001 : AO2 port map( A => v_RAM_OUT0_23_port, B => n1675, C => n4922, D => 
                           n4578, Z => n1671);
   U5002 : AO3 port map( A => n1646, B => n1667, C => n1668, D => n1669, Z => 
                           n4233);
   U5003 : AO7 port map( A => v_KEY_COLUMN_19_port, B => n1609, C => n1650, Z 
                           => n1670);
   U5004 : AO3 port map( A => n1646, B => n1661, C => n1662, D => n1663, Z => 
                           n4234);
   U5005 : AO7 port map( A => n4664, B => n1609, C => n1650, Z => n1666);
   U5006 : AO3 port map( A => n4903, B => n1646, C => n1658, D => n1659, Z => 
                           n4235);
   U5007 : AO7 port map( A => v_KEY_COLUMN_21_port, B => n1609, C => n1650, Z 
                           => n1660);
   U5008 : AO3 port map( A => n1646, B => n1651, C => n1652, D => n1653, Z => 
                           n4236);
   U5009 : AO7 port map( A => n4665, B => n1609, C => n1650, Z => n1656);
   U5010 : AO3 port map( A => n1645, B => n1646, C => n1647, D => n1648, Z => 
                           n4237);
   U5011 : AO7 port map( A => n4666, B => n1609, C => n1650, Z => n1649);
   U5012 : AO3 port map( A => n1553, B => n1726, C => n1748, D => n1749, Z => 
                           n4239);
   U5013 : AO7 port map( A => v_KEY_COLUMN_9_port, B => n1609, C => n1731, Z =>
                           n1750);
   U5014 : AO3 port map( A => n1549, B => n1726, C => n1745, D => n1746, Z => 
                           n4240);
   U5015 : AO7 port map( A => n4658, B => n1609, C => n1731, Z => n1747);
   U5016 : AO3 port map( A => n1544, B => n1726, C => n1742, D => n1743, Z => 
                           n4241);
   U5017 : AO7 port map( A => n4659, B => n1609, C => n1731, Z => n1744);
   U5018 : AO3 port map( A => n1540, B => n1726, C => n1739, D => n1740, Z => 
                           n4242);
   U5019 : AO7 port map( A => v_KEY_COLUMN_12_port, B => n1609, C => n1731, Z 
                           => n1741);
   U5020 : AO3 port map( A => n1535, B => n1726, C => n1735, D => n1736, Z => 
                           n4243);
   U5021 : AO7 port map( A => n4660, B => n1609, C => n1731, Z => n1738);
   U5022 : AO3 port map( A => n1530, B => n1726, C => n1732, D => n1733, Z => 
                           n4244);
   U5023 : AO7 port map( A => n4661, B => n1609, C => n1731, Z => n1734);
   U5024 : AO3 port map( A => n1522, B => n1726, C => n1727, D => n1728, Z => 
                           n4245);
   U5025 : AO7 port map( A => n4662, B => n1609, C => n1731, Z => n1730);
   U5026 : AO3 port map( A => n1598, B => n1755, C => n1780, D => n1781, Z => 
                           n4246);
   U5027 : AO7 port map( A => v_KEY_COLUMN_0_port, B => n1609, C => n1759, Z =>
                           n1782);
   U5028 : AO3 port map( A => n1589, B => n1755, C => n1773, D => n1774, Z => 
                           n4248);
   U5029 : AO7 port map( A => v_KEY_COLUMN_2_port, B => n1609, C => n1759, Z =>
                           n1775);
   U5030 : AO3 port map( A => n1585, B => n1755, C => n1770, D => n1771, Z => 
                           n4249);
   U5031 : AO7 port map( A => v_KEY_COLUMN_3_port, B => n1609, C => n1759, Z =>
                           n1772);
   U5032 : AO3 port map( A => n1581, B => n1755, C => n1767, D => n1768, Z => 
                           n4250);
   U5033 : AO7 port map( A => v_KEY_COLUMN_4_port, B => n1609, C => n1759, Z =>
                           n1769);
   U5034 : AO3 port map( A => n1570, B => n1755, C => n1760, D => n1761, Z => 
                           n4252);
   U5035 : AO7 port map( A => n4656, B => n1609, C => n1759, Z => n1762);
   U5036 : AO3 port map( A => n1563, B => n1755, C => n1756, D => n1757, Z => 
                           n4253);
   U5037 : AO7 port map( A => n4657, B => n1609, C => n1759, Z => n1758);
   U5038 : AO3 port map( A => n1640, B => n1783, C => n1808, D => n1809, Z => 
                           n4254);
   U5039 : AO7 port map( A => n4667, B => n4352, C => n1788, Z => n1810);
   U5040 : AO3 port map( A => n1636, B => n1783, C => n1805, D => n1806, Z => 
                           n4255);
   U5041 : AO7 port map( A => v_KEY_COLUMN_25_port, B => n4352, C => n1788, Z 
                           => n1807);
   U5042 : AO3 port map( A => n1612, B => n1783, C => n1789, D => n1790, Z => 
                           n4260);
   U5043 : AO7 port map( A => n4670, B => n4352, C => n1788, Z => n1791);
   U5044 : AO3 port map( A => n1811, B => n1837, C => n1838, D => n1839, Z => 
                           n4262);
   U5045 : AO7 port map( A => v_KEY_COLUMN_16_port, B => n4352, C => n1815, Z 
                           => n1840);
   U5046 : AO3 port map( A => n1694, B => n1811, C => n1834, D => n1835, Z => 
                           n4263);
   U5047 : AO7 port map( A => n4663, B => n4352, C => n1815, Z => n1836);
   U5048 : AO3 port map( A => n1645, B => n1811, C => n1812, D => n1813, Z => 
                           n4269);
   U5049 : AO7 port map( A => n4666, B => n4352, C => n1815, Z => n1814);
   U5050 : AO3 port map( A => n1553, B => n1841, C => n1882, D => n1883, Z => 
                           n4271);
   U5051 : AO7 port map( A => v_KEY_COLUMN_9_port, B => n4352, C => n1846, Z =>
                           n1885);
   U5052 : AO3 port map( A => n1860, B => n1841, C => n1861, D => n1862, Z => 
                           n4272);
   U5053 : AO6 port map( A => n4905, B => v_RAM_OUT0_9_port, C => n1865, Z => 
                           n1860);
   U5054 : AO3 port map( A => n1544, B => n1841, C => n1857, D => n1858, Z => 
                           n4273);
   U5055 : AO7 port map( A => n4659, B => n4352, C => n1846, Z => n1859);
   U5056 : AO3 port map( A => n1540, B => n1841, C => n1854, D => n1855, Z => 
                           n4274);
   U5057 : AO7 port map( A => v_KEY_COLUMN_12_port, B => n4352, C => n1846, Z 
                           => n1856);
   U5058 : AO3 port map( A => n1535, B => n1841, C => n1850, D => n1851, Z => 
                           n4275);
   U5059 : AO7 port map( A => n4660, B => n4352, C => n1846, Z => n1853);
   U5060 : AO3 port map( A => n1530, B => n1841, C => n1847, D => n1848, Z => 
                           n4276);
   U5061 : AO7 port map( A => n4661, B => n4352, C => n1846, Z => n1849);
   U5062 : AO3 port map( A => n1522, B => n1841, C => n1842, D => n1843, Z => 
                           n4277);
   U5063 : AO7 port map( A => n4662, B => n4352, C => n1846, Z => n1845);
   U5064 : AO3 port map( A => n1598, B => n3295, C => n3668, D => n3669, Z => 
                           n4278);
   U5065 : AO7 port map( A => v_KEY_COLUMN_0_port, B => n4352, C => n3299, Z =>
                           n3670);
   U5066 : AO3 port map( A => n1593, B => n3295, C => n3629, D => n3630, Z => 
                           n4279);
   U5067 : AO7 port map( A => v_KEY_COLUMN_1_port, B => n4352, C => n3299, Z =>
                           n3632);
   U5068 : AO3 port map( A => n1570, B => n3295, C => n3373, D => n3374, Z => 
                           n4284);
   U5069 : AO7 port map( A => n4656, B => n4352, C => n3299, Z => n3375);
   U5070 : AO3 port map( A => n1563, B => n3295, C => n3296, D => n3297, Z => 
                           n4285);
   U5071 : AO7 port map( A => n4657, B => n4352, C => n3299, Z => n3298);
   U5072 : NR3 port map( A => n1459, B => n4849, C => n4852, Z => n1450);
   U5073 : AO7 port map( A => v_RAM_OUT0_31_port, B => n2746, C => n2747, Z => 
                           n1627);
   U5074 : AO6 port map( A => v_RAM_OUT0_29_port, B => n2769, C => n2770, Z => 
                           n2746);
   U5075 : AO3 port map( A => n2748, B => n2749, C => v_RAM_OUT0_31_port, D => 
                           n2750, Z => n2747);
   U5076 : AO4 port map( A => n2771, B => n4689, C => n2772, D => n4688, Z => 
                           n2770);
   U5077 : AO7 port map( A => v_RAM_OUT0_23_port, B => n3150, C => n3151, Z => 
                           n1667);
   U5078 : AO6 port map( A => v_RAM_OUT0_21_port, B => n3173, C => n3174, Z => 
                           n3150);
   U5079 : AO3 port map( A => n3152, B => n3153, C => v_RAM_OUT0_23_port, D => 
                           n3154, Z => n3151);
   U5080 : AO4 port map( A => n3175, B => n4684, C => n3176, D => n4685, Z => 
                           n3174);
   U5081 : AO7 port map( A => v_RAM_OUT0_7_port, B => n3551, C => n3552, Z => 
                           n1585);
   U5082 : AO6 port map( A => v_RAM_OUT0_5_port, B => n3574, C => n3575, Z => 
                           n3551);
   U5083 : AO3 port map( A => n3553, B => n3554, C => v_RAM_OUT0_7_port, D => 
                           n3555, Z => n3552);
   U5084 : AO4 port map( A => n3576, B => n4680, C => n3577, D => n4681, Z => 
                           n3575);
   U5085 : AO4 port map( A => v_RAM_OUT0_31_port, B => n4867, C => n1942, D => 
                           n4587, Z => n1632);
   U5086 : AO6 port map( A => v_RAM_OUT0_29_port, B => n1944, C => n1945, Z => 
                           n1942);
   U5087 : AO4 port map( A => n4865, B => n4688, C => n1948, D => n4689, Z => 
                           n1945);
   U5088 : AO4 port map( A => v_RAM_OUT0_23_port, B => n4922, C => n3195, D => 
                           n4578, Z => n1830);
   U5089 : AO6 port map( A => v_RAM_OUT0_21_port, B => n1679, C => n3196, Z => 
                           n3195);
   U5090 : AO4 port map( A => n4930, B => n4685, C => n3197, D => n4684, Z => 
                           n3196);
   U5091 : AO4 port map( A => v_RAM_OUT0_7_port, B => n5004, C => n3596, D => 
                           n4588, Z => n1589);
   U5092 : AO6 port map( A => v_RAM_OUT0_5_port, B => n2445, C => n3597, Z => 
                           n3596);
   U5093 : AO4 port map( A => n5012, B => n4681, C => n3598, D => n4680, Z => 
                           n3597);
   U5094 : NR4 port map( A => n1893, B => n1894, C => n4569, D => n1895, Z => 
                           n1892);
   U5095 : AO4 port map( A => n1896, B => n1897, C => n4691, D => n1899, Z => 
                           n1894);
   U5096 : AO2 port map( A => n1910, B => n4378, C => v_RAM_OUT0_10_port, D => 
                           n1911, Z => n1909);
   U5097 : AO4 port map( A => n2403, B => n2074, C => n1912, D => n2404, Z => 
                           n1895);
   U5098 : AO7 port map( A => n2407, B => n4707, C => n2087_port, Z => n2406);
   U5099 : IVDA port map( A => n1973, Y => n4511, Z => n4686);
   U5100 : AO4 port map( A => n2640, B => n2641, C => v_RAM_OUT0_31_port, D => 
                           n2642, Z => n2639);
   U5101 : AO6 port map( A => n2522, B => n2584, C => n5059, Z => n2783);
   U5102 : AO6 port map( A => n2926, B => n2987, C => n5056, Z => n3188);
   U5103 : AO6 port map( A => n3328, B => n3388, C => n5050, Z => n3589);
   U5104 : AO7 port map( A => n1906, B => n4359, C => n2110, Z => n2243);
   U5105 : AO3 port map( A => n2245, B => n4707, C => n2246, D => n4906, Z => 
                           n2244);
   U5106 : AO2 port map( A => n4701, B => n4955, C => n4360, D => n4970, Z => 
                           n2246);
   U5107 : AO2 port map( A => n2667, B => n4686, C => n4900, D => 
                           v_RAM_OUT0_28_port, Z => n2666);
   U5108 : AO4 port map( A => n4892, B => n4687, C => n4902, D => n2513, Z => 
                           n2510);
   U5109 : AO6 port map( A => n4896, B => v_RAM_OUT0_26_port, C => n4371, Z => 
                           n2513);
   U5110 : AO4 port map( A => n4917, B => n4682, C => n4927, D => n2917, Z => 
                           n2914);
   U5111 : AO6 port map( A => n4934, B => v_RAM_OUT0_18_port, C => n4369, Z => 
                           n2917);
   U5112 : AO4 port map( A => n4412, B => n4707, C => n4359, D => n4958, Z => 
                           n2369);
   U5113 : AO4 port map( A => v_RAM_OUT0_10_port, B => n2093, C => n4359, D => 
                           n2094, Z => n2091);
   U5114 : AO4 port map( A => n4999, B => n4678, C => n5009, D => n3319, Z => 
                           n3316);
   U5115 : AO6 port map( A => n5016, B => v_RAM_OUT0_2_port, C => n4370, Z => 
                           n3319);
   U5116 : EO1 port map( A => n4412, B => n4360, C => n2234, D => n4359, Z => 
                           n2421);
   U5117 : AO6 port map( A => n1902, B => n4378, C => n1904, Z => n1896);
   U5118 : EON1 port map( A => n4707, B => n1906, C => n1907, D => n4360, Z => 
                           n1904);
   U5119 : AO2 port map( A => n4906, B => n2337, C => n2338, D => n2339, Z => 
                           n2336);
   U5120 : AO3 port map( A => n2215, B => n4361, C => n2341, D => n2343, Z => 
                           n2337);
   U5121 : AO2 port map( A => n5040, B => n2332, C => n1876, D => n5039, Z => 
                           n2327);
   U5122 : AO6 port map( A => n1870, B => v_RAM_OUT0_13_port, C => n2294, Z => 
                           n2328);
   U5123 : AO3 port map( A => n4411, B => n2519, C => n2840, D => n2841, Z => 
                           n2829);
   U5124 : AO2 port map( A => n5060, B => n2523, C => n4878, D => n5061, Z => 
                           n2841);
   U5125 : AO2 port map( A => n2842, B => n2531, C => n4901, D => n2527, Z => 
                           n2840);
   U5126 : AO3 port map( A => n4914, B => n2585, C => v_RAM_OUT0_29_port, D => 
                           n2838, Z => n2830);
   U5127 : EO1 port map( A => n2655, B => n2522, C => n2530, D => n1958, Z => 
                           n2838);
   U5128 : AO7 port map( A => n2628, B => n2629, C => n5042, Z => n2627);
   U5129 : AO3 port map( A => n4866, B => n1959, C => n2630, D => n2625, Z => 
                           n2628);
   U5130 : AO4 port map( A => n1977, B => n4704, C => v_RAM_OUT0_28_port, D => 
                           n2562, Z => n2629);
   U5131 : AO3 port map( A => n4406, B => n2923, C => n3244, D => n3245, Z => 
                           n3233);
   U5132 : AO2 port map( A => n5057, B => n2927, C => n4940, D => n5053, Z => 
                           n3245);
   U5133 : AO2 port map( A => n3246, B => n2938, C => n4926, D => n2932, Z => 
                           n3244);
   U5134 : AO3 port map( A => n4925, B => n2988, C => v_RAM_OUT0_21_port, D => 
                           n3242, Z => n3234);
   U5135 : EO1 port map( A => n3060, B => n2926, C => n2936, D => n1689, Z => 
                           n3242);
   U5136 : AO2 port map( A => n4989, B => v_RAM_OUT0_10_port, C => n2065, D => 
                           n2276, Z => n2275);
   U5137 : AO6 port map( A => n2176, B => n2177, C => n1897, Z => n2175);
   U5138 : EO1 port map( A => n4701, B => n2178, C => n2179, D => 
                           v_RAM_OUT0_10_port, Z => n2177);
   U5139 : AO2 port map( A => n4956, B => n4360, C => n4379, D => n2047, Z => 
                           n2176);
   U5140 : AO3 port map( A => n4405, B => n3325, C => n3646, D => n3647, Z => 
                           n3635);
   U5141 : AO2 port map( A => n5051, B => n3329, C => n5022, D => n5047, Z => 
                           n3647);
   U5142 : AO2 port map( A => n3648, B => n3340, C => n5008, D => n3334, Z => 
                           n3646);
   U5143 : AO3 port map( A => n5007, B => n3389, C => v_RAM_OUT0_5_port, D => 
                           n3644, Z => n3636);
   U5144 : EO1 port map( A => n3462, B => n3328, C => n3338, D => n2455, Z => 
                           n3644);
   U5145 : AO7 port map( A => n3433, B => n3434, C => n5044, Z => n3432);
   U5146 : AO3 port map( A => n5027, B => n3359, C => n3435, D => n3429, Z => 
                           n3433);
   U5147 : AO4 port map( A => n2489, B => n4695, C => v_RAM_OUT0_4_port, D => 
                           n3367, Z => n3434);
   U5148 : AO7 port map( A => n4408, B => n2469, C => n2470, Z => n2468);
   U5149 : AO2 port map( A => n4505, B => n2471, C => n5006, D => n4400, Z => 
                           n2470);
   U5150 : AO4 port map( A => n5046, B => n2474, C => n2475, D => n2476, Z => 
                           n2471);
   U5151 : AO2 port map( A => v_RAM_OUT0_2_port, B => n2477, C => n5000, D => 
                           n4363, Z => n2475);
   U5152 : AO7 port map( A => v_RAM_OUT0_5_port, B => n2480, C => n2481, Z => 
                           n2467);
   U5153 : AO2 port map( A => n5045, B => n2483, C => n2484, D => n5044, Z => 
                           n2481);
   U5154 : AO4 port map( A => n5046, B => n2486, C => n2487, D => n2476, Z => 
                           n2483);
   U5155 : AO2 port map( A => v_RAM_OUT0_2_port, B => n4679, C => n2489, D => 
                           n4363, Z => n2487);
   U5156 : AO7 port map( A => n4410, B => n1982, C => n2869, Z => n2868);
   U5157 : AO2 port map( A => n4503, B => n2870, C => n4874, D => n4399, Z => 
                           n2869);
   U5158 : AO4 port map( A => n5058, B => n1986, C => n2876, D => n1978, Z => 
                           n2870);
   U5159 : AO2 port map( A => v_RAM_OUT0_26_port, B => n1988, C => n4885, D => 
                           n4362, Z => n2876);
   U5160 : AO7 port map( A => v_RAM_OUT0_29_port, B => n1970, C => n2884, Z => 
                           n2867);
   U5161 : AO2 port map( A => n5043, B => n2885, C => n1980, D => n5042, Z => 
                           n2884);
   U5162 : AO4 port map( A => n5058, B => n2540, C => n2888, D => n1978, Z => 
                           n2885);
   U5163 : AO2 port map( A => v_RAM_OUT0_26_port, B => n4686, C => n1977, D => 
                           n4362, Z => n2888);
   U5164 : AO7 port map( A => n4409, B => n1705, C => n1706, Z => n1704);
   U5165 : AO2 port map( A => n4504, B => n1707, C => n4924, D => n4402, Z => 
                           n1706);
   U5166 : AO4 port map( A => n5052, B => n1710, C => n1711, D => n1712, Z => 
                           n1707);
   U5167 : AO2 port map( A => v_RAM_OUT0_18_port, B => n1713, C => n4918, D => 
                           n4365, Z => n1711);
   U5168 : AO7 port map( A => v_RAM_OUT0_21_port, B => n1716, C => n1717, Z => 
                           n1703);
   U5169 : AO2 port map( A => n5038, B => n1719, C => n1720, D => n5037, Z => 
                           n1717);
   U5170 : AO4 port map( A => n5052, B => n1722, C => n1723, D => n1712, Z => 
                           n1719);
   U5171 : AO2 port map( A => v_RAM_OUT0_18_port, B => n4683, C => n1725, D => 
                           n4365, Z => n1723);
   U5172 : AO6 port map( A => n2658, B => n2659, C => n4410, Z => n2643);
   U5173 : AO2 port map( A => v_RAM_OUT0_25_port, B => n2663, C => n4891, D => 
                           n5063, Z => n2658);
   U5174 : AO3 port map( A => n1977, B => n4705, C => n2660, D => n2661, Z => 
                           n2659);
   U5175 : AO4 port map( A => n4362, B => n2665, C => v_RAM_OUT0_26_port, D => 
                           n2666, Z => n2663);
   U5176 : AO3 port map( A => n4700, B => n3022, C => n4402, D => n3023, Z => 
                           n3012);
   U5177 : AO6 port map( A => n3027, B => n3028, C => n4682, Z => n3026);
   U5178 : AO3 port map( A => v_RAM_OUT0_8_port, B => n2110, C => n2111, D => 
                           n2112, Z => n2109);
   U5179 : AO2 port map( A => n2113, B => n4379, C => n4955, D => n4701, Z => 
                           n2112);
   U5180 : AO2 port map( A => n2114, B => n4360, C => n4993, D => n4702, Z => 
                           n2111);
   U5181 : AO3 port map( A => n1632, B => n1783, C => n1802, D => n1803, Z => 
                           n4256);
   U5182 : AO7 port map( A => v_KEY_COLUMN_26_port, B => n4352, C => n1788, Z 
                           => n1804);
   U5183 : AO3 port map( A => n1627, B => n1783, C => n1799, D => n1800, Z => 
                           n4257);
   U5184 : AO7 port map( A => n4668, B => n4352, C => n1788, Z => n1801);
   U5185 : AO3 port map( A => n4870, B => n1783, C => n1792, D => n1793, Z => 
                           n4259);
   U5186 : AO7 port map( A => v_KEY_COLUMN_29_port, B => n4352, C => n1788, Z 
                           => n1794);
   U5187 : AO3 port map( A => n1811, B => n1830, C => n1831, D => n1832, Z => 
                           n4264);
   U5188 : AO7 port map( A => v_KEY_COLUMN_18_port, B => n4352, C => n1815, Z 
                           => n1833);
   U5189 : AO3 port map( A => n1667, B => n1811, C => n1827, D => n1828, Z => 
                           n4265);
   U5190 : AO7 port map( A => v_KEY_COLUMN_19_port, B => n4352, C => n1815, Z 
                           => n1829);
   U5191 : AO3 port map( A => n4903, B => n1811, C => n1820, D => n1821, Z => 
                           n4267);
   U5192 : AO7 port map( A => v_KEY_COLUMN_21_port, B => n4352, C => n1815, Z 
                           => n1822);
   U5193 : AO3 port map( A => n1589, B => n3295, C => n3593, D => n3594, Z => 
                           n4280);
   U5194 : AO7 port map( A => v_KEY_COLUMN_2_port, B => n4352, C => n3299, Z =>
                           n3595);
   U5195 : AO3 port map( A => n1585, B => n3295, C => n3548, D => n3549, Z => 
                           n4281);
   U5196 : AO7 port map( A => v_KEY_COLUMN_3_port, B => n4352, C => n3299, Z =>
                           n3550);
   U5197 : AO3 port map( A => n1581, B => n3295, C => n3502, D => n3503, Z => 
                           n4282);
   U5198 : AO7 port map( A => v_KEY_COLUMN_4_port, B => n4352, C => n3299, Z =>
                           n3504);
   U5199 : AO3 port map( A => n4911, B => n3295, C => n3441, D => n3442, Z => 
                           n4283);
   U5200 : AO7 port map( A => n4655, B => n4352, C => n3299, Z => n3444);
   U5201 : ND4 port map( A => n2996, B => n2997, C => n2998, D => n2999, Z => 
                           n2978);
   U5202 : AO2 port map( A => n4951, B => n5054, C => n5057, D => n3007, Z => 
                           n2998);
   U5203 : AO2 port map( A => n5055, B => n3011, C => n2968, D => n5056, Z => 
                           n2996);
   U5204 : AO2 port map( A => n3000, B => v_RAM_OUT0_17_port, C => n4945, D => 
                           n4498, Z => n2999);
   U5205 : ND4 port map( A => n2050, B => v_RAM_OUT0_15_port, C => n2051, D => 
                           n2052, Z => n2027);
   U5206 : AO2 port map( A => n2065, B => n2066, C => n5041, D => n2067, Z => 
                           n2050);
   U5207 : AO2 port map( A => n2054, B => n1914, C => v_RAM_OUT0_13_port, D => 
                           n2055, Z => n2051);
   U5208 : ND4 port map( A => n2722, B => n2723, C => n2724, D => n2725, Z => 
                           n2699);
   U5209 : ND4 port map( A => n2701, B => v_RAM_OUT0_31_port, C => n2702, D => 
                           n2703, Z => n2700);
   U5210 : AO7 port map( A => n2726, B => n2727, C => n5043, Z => n2725);
   U5211 : ND4 port map( A => n3126, B => n3127, C => n3128, D => n3129, Z => 
                           n3104);
   U5212 : ND4 port map( A => n3106, B => v_RAM_OUT0_23_port, C => n3107, D => 
                           n3108, Z => n3105);
   U5213 : AO7 port map( A => n3130, B => n3131, C => n5038, Z => n3129);
   U5214 : ND4 port map( A => n3527, B => n3528, C => n3529, D => n3530, Z => 
                           n3505);
   U5215 : ND4 port map( A => n3507, B => v_RAM_OUT0_7_port, C => n3508, D => 
                           n3509, Z => n3506);
   U5216 : AO7 port map( A => n3531, B => n3532, C => n5045, Z => n3530);
   U5217 : AO4 port map( A => n4689, B => n2552, C => n4688, D => n4686, Z => 
                           n2547);
   U5218 : AO4 port map( A => n4684, B => n2955, C => n4685, D => n4683, Z => 
                           n2951);
   U5219 : AO4 port map( A => n4680, B => n3357, C => n4681, D => n4679, Z => 
                           n3353);
   U5220 : ND4 port map( A => n2889, B => n2890, C => n2891, D => n2892, Z => 
                           n1970);
   U5221 : AO2 port map( A => n5060, B => n4411, C => n5059, D => n2822, Z => 
                           n2889);
   U5222 : AO2 port map( A => n4914, B => n5062, C => n2531, D => n2618, Z => 
                           n2892);
   U5223 : ND4 port map( A => n3273, B => n3274, C => n3275, D => n3276, Z => 
                           n1716);
   U5224 : AO2 port map( A => n5057, B => n4406, C => n5056, D => n3208, Z => 
                           n3273);
   U5225 : AO2 port map( A => n4925, B => n5054, C => n2938, D => n3020, Z => 
                           n3276);
   U5226 : ND4 port map( A => n3677, B => n3678, C => n3679, D => n3680, Z => 
                           n2480);
   U5227 : AO2 port map( A => n5051, B => n4405, C => n5050, D => n3609, Z => 
                           n3677);
   U5228 : AO2 port map( A => n5007, B => n5048, C => n3340, D => n3421, Z => 
                           n3680);
   U5229 : EON1 port map( A => v_RAM_OUT0_10_port, B => n2130, C => n4702, D =>
                           n2061, Z => n2126);
   U5230 : AO3 port map( A => n4707, B => n2056, C => n2057, D => n2058, Z => 
                           n2055);
   U5231 : AO2 port map( A => n4702, B => n2060, C => n2061, D => n4404, Z => 
                           n2058);
   U5232 : NR3 port map( A => n4883, B => n2886, C => n2887, Z => n1980);
   U5233 : AO4 port map( A => n1959, B => n4686, C => n4894, D => n4705, Z => 
                           n2886);
   U5234 : AO4 port map( A => v_RAM_OUT0_28_port, B => n2528, C => n2652, D => 
                           n4687, Z => n2887);
   U5235 : NR3 port map( A => n5065, B => n3279, C => n3280, Z => n1720);
   U5236 : AO4 port map( A => n2957, B => n4683, C => n4951, D => n4700, Z => 
                           n3279);
   U5237 : AO4 port map( A => v_RAM_OUT0_20_port, B => n2933, C => n3056, D => 
                           n4682, Z => n3280);
   U5238 : NR3 port map( A => n5070, B => n3683, C => n3684, Z => n2484);
   U5239 : AO4 port map( A => n3359, B => n4679, C => n5033, D => n4697, Z => 
                           n3683);
   U5240 : AO4 port map( A => v_RAM_OUT0_4_port, B => n3335, C => n3458, D => 
                           n4678, Z => n3684);
   U5241 : AO3 port map( A => n2759, B => n2651, C => v_RAM_OUT0_29_port, D => 
                           n2760, Z => n2749);
   U5242 : AO2 port map( A => n5062, B => n2568, C => n2522, D => n2761, Z => 
                           n2760);
   U5243 : AO2 port map( A => n5042, B => n2716, C => n4399, D => n2717, Z => 
                           n2701);
   U5244 : AO3 port map( A => v_RAM_OUT0_26_port, B => n2562, C => n4875, D => 
                           n2720, Z => n2716);
   U5245 : AO3 port map( A => n4704, B => n2706, C => n1959, D => n2718, Z => 
                           n2717);
   U5246 : AO2 port map( A => n4882, B => n4357, C => n4371, D => n2721, Z => 
                           n2720);
   U5247 : AO3 port map( A => n3163, B => n3055, C => v_RAM_OUT0_21_port, D => 
                           n3164, Z => n3153);
   U5248 : AO2 port map( A => n5054, B => n2970, C => n2926, D => n3165, Z => 
                           n3164);
   U5249 : AO2 port map( A => n5037, B => n3120, C => n4402, D => n3121, Z => 
                           n3106);
   U5250 : AO3 port map( A => v_RAM_OUT0_18_port, B => n2965, C => n4931, D => 
                           n3124, Z => n3120);
   U5251 : AO3 port map( A => n4698, B => n3111, C => n2957, D => n3122, Z => 
                           n3121);
   U5252 : AO2 port map( A => n4954, B => n4355, C => n4369, D => n3125, Z => 
                           n3124);
   U5253 : AO7 port map( A => n2288, B => n2289, C => v_RAM_OUT0_13_port, Z => 
                           n2287);
   U5254 : AO4 port map( A => n4994, B => n4690, C => n2291, D => n4361, Z => 
                           n2288);
   U5255 : AO4 port map( A => n2066, B => n4707, C => n4359, D => n2290, Z => 
                           n2289);
   U5256 : AO3 port map( A => n3564, B => n3457, C => v_RAM_OUT0_5_port, D => 
                           n3565, Z => n3554);
   U5257 : AO2 port map( A => n5048, B => n3372, C => n3328, D => n3566, Z => 
                           n3565);
   U5258 : AO2 port map( A => n5044, B => n3521, C => n4400, D => n3522, Z => 
                           n3507);
   U5259 : AO3 port map( A => v_RAM_OUT0_2_port, B => n3367, C => n5013, D => 
                           n3525, Z => n3521);
   U5260 : AO3 port map( A => n4695, B => n3512, C => n3359, D => n3523, Z => 
                           n3522);
   U5261 : AO2 port map( A => n5036, B => n4356, C => n4370, D => n3526, Z => 
                           n3525);
   U5262 : AO7 port map( A => n4408, B => n2445, C => n2446, Z => n2441);
   U5263 : AO2 port map( A => n5012, B => n4505, C => n4400, D => n2450, Z => 
                           n2446);
   U5264 : AO2 port map( A => n5024, B => n4373, C => n5035, D => 
                           v_RAM_OUT0_2_port, Z => n2451);
   U5265 : AO7 port map( A => n4410, B => n1944, C => n2809, Z => n2791);
   U5266 : AO2 port map( A => n4865, B => n4503, C => n4399, D => n2810, Z => 
                           n2809);
   U5267 : AO2 port map( A => n4881, B => n4372, C => n4898, D => 
                           v_RAM_OUT0_26_port, Z => n2811);
   U5268 : AO7 port map( A => n4409, B => n1679, C => n1680, Z => n1675);
   U5269 : AO2 port map( A => n4930, B => n4504, C => n4402, D => n1684, Z => 
                           n1680);
   U5270 : AO2 port map( A => n4942, B => n4374, C => n4953, D => 
                           v_RAM_OUT0_18_port, Z => n1685);
   U5271 : AO3 port map( A => n1978, B => n2676, C => n2814, D => n2815, Z => 
                           n2813);
   U5272 : AO2 port map( A => n4873, B => n4357, C => n4866, D => n4372, Z => 
                           n2815);
   U5273 : AO3 port map( A => n1712, B => n3081, C => n3201, D => n3202, Z => 
                           n3200);
   U5274 : AO2 port map( A => n4950, B => n4355, C => n4945, D => n4374, Z => 
                           n3202);
   U5275 : AO3 port map( A => n2476, B => n3483, C => n3602, D => n3603, Z => 
                           n3601);
   U5276 : AO2 port map( A => n5032, B => n4356, C => n5027, D => n4373, Z => 
                           n3603);
   U5277 : AO3 port map( A => n4404, B => n2226, C => n2227, D => n2228, Z => 
                           n2225);
   U5278 : AO2 port map( A => n2191, B => n4360, C => n2211, D => n4702, Z => 
                           n2228);
   U5279 : AO3 port map( A => n2032, B => n4378, C => n2033, D => n4707, Z => 
                           n2031);
   U5280 : AO7 port map( A => v_RAM_OUT0_10_port, B => n4981, C => n4359, Z => 
                           n2035);
   U5281 : AO3 port map( A => n4925, B => n4700, C => n4504, D => n3014, Z => 
                           n3013);
   U5282 : AO6 port map( A => n3019, B => n3020, C => n4698, Z => n3017);
   U5283 : EON1 port map( A => n4384, B => n1454, C => N2085, D => n1450, Z => 
                           n4307);
   U5284 : EON1 port map( A => n4601, B => n1454, C => n4601, D => n1450, Z => 
                           n4310);
   U5285 : ND4 port map( A => n2594, B => n2595, C => n2596, D => n2597, Z => 
                           n2576);
   U5286 : AO2 port map( A => n4894, B => n5062, C => n5060, D => n1955, Z => 
                           n2596);
   U5287 : AO2 port map( A => n5063, B => n2608, C => n2565, D => n5059, Z => 
                           n2594);
   U5288 : AO2 port map( A => n2598, B => v_RAM_OUT0_25_port, C => n4866, D => 
                           n4499, Z => n2597);
   U5289 : ND4 port map( A => n3397, B => n3398, C => n3399, D => n3400, Z => 
                           n3379);
   U5290 : AO2 port map( A => n5033, B => n5048, C => n5051, D => n3408, Z => 
                           n3399);
   U5291 : AO2 port map( A => n5049, B => n3412, C => n3370, D => n5050, Z => 
                           n3397);
   U5292 : AO2 port map( A => n3401, B => v_RAM_OUT0_1_port, C => n5027, D => 
                           n4497, Z => n3400);
   U5293 : ND3 port map( A => n3062, B => n4365, C => v_RAM_OUT0_17_port, Z => 
                           n3061);
   U5294 : ND3 port map( A => n3464, B => n4363, C => v_RAM_OUT0_1_port, Z => 
                           n3463);
   U5295 : AO7 port map( A => v_RAM_OUT0_24_port, B => n4705, C => n4687, Z => 
                           n1951);
   U5296 : AO7 port map( A => v_RAM_OUT0_16_port, B => n4700, C => n4682, Z => 
                           n1687);
   U5297 : AO7 port map( A => v_RAM_OUT0_0_port, B => n4697, C => n4678, Z => 
                           n2453);
   U5298 : IVDA port map( A => n1947, Y => n4503, Z => n4688);
   U5299 : IVDA port map( A => n2906, Y => n4504, Z => n4685);
   U5300 : IVDA port map( A => n3308, Y => n4505, Z => n4681);
   U5301 : IVDA port map( A => n1898, Y => n4506, Z => n4691);
   U5302 : AO6 port map( A => n2120, B => n2121, C => n4707, Z => n2119);
   U5303 : AO6 port map( A => n2965, B => n3082, C => n4700, Z => n3079);
   U5304 : AO6 port map( A => n3367, B => n3484, C => n4697, Z => n3481);
   U5305 : AO6 port map( A => n2738, B => n2739, C => n1959, Z => n2736);
   U5306 : AO6 port map( A => n3142, B => n3143, C => n2957, Z => n3140);
   U5307 : AO6 port map( A => n3543, B => n3544, C => n3359, Z => n3541);
   U5308 : AO2 port map( A => n1507, B => n4529, C => n4858, D => n4423, Z => 
                           n3790);
   U5309 : AO2 port map( A => n1506, B => n4553, C => n1508, D => n4454, Z => 
                           n3791);
   U5310 : AO2 port map( A => n1507, B => n4429, C => n4858, D => n4597, Z => 
                           n3779);
   U5311 : AO2 port map( A => n1506, B => n4595, C => n1508, D => n4442, Z => 
                           n3780);
   U5312 : AO2 port map( A => n1507, B => n4430, C => n4858, D => n4533, Z => 
                           n3768);
   U5313 : AO2 port map( A => n1506, B => n4421, C => n1508, D => n4528, Z => 
                           n3769);
   U5314 : AO2 port map( A => n1507, B => n4401, C => n4858, D => n4448, Z => 
                           n3757);
   U5315 : AO2 port map( A => n1506, B => n4554, C => n1508, D => n4443, Z => 
                           n3758);
   U5316 : AO2 port map( A => n1507, B => n4566, C => n4858, D => n4449, Z => 
                           n3746);
   U5317 : AO2 port map( A => n1506, B => n4447, C => n1508, D => n4592, Z => 
                           n3747);
   U5318 : AO2 port map( A => n1507, B => n4414, C => n4858, D => n4598, Z => 
                           n3735);
   U5319 : AO2 port map( A => n1506, B => n4596, C => n1508, D => n4413, Z => 
                           n3736);
   U5320 : AO2 port map( A => n1507, B => n4398, C => n4858, D => n4434, Z => 
                           n3724);
   U5321 : AO2 port map( A => n1506, B => n4397, C => n1508, D => n4428, Z => 
                           n3725);
   U5322 : AO2 port map( A => n1507, B => n4418, C => n4858, D => n4599, Z => 
                           n3712);
   U5323 : AO2 port map( A => n1506, B => n4422, C => n1508, D => n4593, Z => 
                           n3713);
   U5324 : AO6 port map( A => n5042, B => n2730, C => v_RAM_OUT0_31_port, Z => 
                           n2724);
   U5325 : AO3 port map( A => n4704, B => n2549, C => n2731, D => n2732, Z => 
                           n2730);
   U5326 : AO7 port map( A => n4887, B => n4897, C => n4703, Z => n2731);
   U5327 : AO2 port map( A => n4902, B => n4357, C => n4371, D => n2619, Z => 
                           n2732);
   U5328 : AO3 port map( A => n4705, B => n2654, C => n4503, D => n2734, Z => 
                           n2723);
   U5329 : AO6 port map( A => n2584, B => n2583, C => n4704, Z => n2737);
   U5330 : AO6 port map( A => n5037, B => n3134, C => v_RAM_OUT0_23_port, Z => 
                           n3128);
   U5331 : AO3 port map( A => n4698, B => n2953, C => n3135, D => n3136, Z => 
                           n3134);
   U5332 : AO7 port map( A => n4928, B => n5066, C => n4699, Z => n3135);
   U5333 : AO2 port map( A => n4927, B => n4355, C => n4369, D => n3022, Z => 
                           n3136);
   U5334 : AO3 port map( A => n4700, B => n3058, C => n4504, D => n3138, Z => 
                           n3127);
   U5335 : AO6 port map( A => n2987, B => n2986, C => n4698, Z => n3141);
   U5336 : AO6 port map( A => n5044, B => n3535, C => v_RAM_OUT0_7_port, Z => 
                           n3529);
   U5337 : AO3 port map( A => n4695, B => n3355, C => n3536, D => n3537, Z => 
                           n3535);
   U5338 : AO7 port map( A => n5010, B => n5071, C => n4696, Z => n3536);
   U5339 : AO2 port map( A => n5009, B => n4356, C => n4370, D => n3423, Z => 
                           n3537);
   U5340 : AO3 port map( A => n4697, B => n3460, C => n4505, D => n3539, Z => 
                           n3528);
   U5341 : AO6 port map( A => n3388, B => n3387, C => n4695, Z => n3542);
   U5342 : AO3 port map( A => n4914, B => n4705, C => n4503, D => n2612, Z => 
                           n2610);
   U5343 : AO6 port map( A => n2617, B => n2618, C => n4704, Z => n2615);
   U5344 : AO3 port map( A => n4705, B => n2619, C => n4399, D => n2620, Z => 
                           n2609);
   U5345 : AO6 port map( A => n2624, B => n2625, C => n4687, Z => n2623);
   U5346 : AO3 port map( A => n5007, B => n4697, C => n4505, D => n3415, Z => 
                           n3414);
   U5347 : AO6 port map( A => n3420, B => n3421, C => n4695, Z => n3418);
   U5348 : AO3 port map( A => n4697, B => n3423, C => n4400, D => n3424, Z => 
                           n3413);
   U5349 : AO6 port map( A => n3428, B => n3429, C => n4678, Z => n3427);
   U5350 : ND3 port map( A => n2657, B => n4362, C => v_RAM_OUT0_25_port, Z => 
                           n2656);
   U5351 : AO6 port map( A => n2562, B => n2677, C => n4705, Z => n2674);
   U5352 : AO4 port map( A => n4687, B => n2617, C => n2729, D => n4705, Z => 
                           n2726);
   U5353 : AO4 port map( A => n4682, B => n3019, C => n3133, D => n4700, Z => 
                           n3130);
   U5354 : AO4 port map( A => n4678, B => n3420, C => n3534, D => n4697, Z => 
                           n3531);
   U5355 : AO2 port map( A => n2709, B => n2689, C => n4503, D => n2710, Z => 
                           n2702);
   U5356 : AO4 port map( A => n4705, B => n2684, C => n4898, D => n2712, Z => 
                           n2710);
   U5357 : AO6 port map( A => n4871, B => v_RAM_OUT0_28_port, C => n4357, Z => 
                           n2712);
   U5358 : AO2 port map( A => n3114, B => n3094, C => n4504, D => n3115, Z => 
                           n3107);
   U5359 : AO4 port map( A => n4700, B => n3089, C => n4953, D => n3116, Z => 
                           n3115);
   U5360 : AO6 port map( A => n4947, B => v_RAM_OUT0_20_port, C => n4355, Z => 
                           n3116);
   U5361 : AO2 port map( A => n3515, B => n3496, C => n4505, D => n3516, Z => 
                           n3508);
   U5362 : AO4 port map( A => n4697, B => n3491, C => n5035, D => n3517, Z => 
                           n3516);
   U5363 : AO6 port map( A => n5029, B => v_RAM_OUT0_4_port, C => n4356, Z => 
                           n3517);
   U5364 : AO4 port map( A => n4464, B => n4349, C => n4710, D => n4621, Z => 
                           n3967);
   U5365 : AO4 port map( A => n4465, B => n4349, C => n4710, D => n4622, Z => 
                           n3973);
   U5366 : AO4 port map( A => n4466, B => n4349, C => n4710, D => n4623, Z => 
                           n3979);
   U5367 : AO4 port map( A => n4467, B => n4349, C => n4710, D => n4624, Z => 
                           n3985);
   U5368 : AO4 port map( A => n4468, B => n4349, C => n4710, D => n4625, Z => 
                           n3991);
   U5369 : AO4 port map( A => n4469, B => n4349, C => n4710, D => n4626, Z => 
                           n3997);
   U5370 : AO4 port map( A => n4470, B => n4349, C => n4710, D => n4627, Z => 
                           n4003);
   U5371 : AO4 port map( A => n4471, B => n4349, C => n4710, D => n4628, Z => 
                           n4009);
   U5372 : AO4 port map( A => n4472, B => n4349, C => n4710, D => n4629, Z => 
                           n4015);
   U5373 : AO4 port map( A => n4473, B => n4349, C => n4710, D => n4630, Z => 
                           n4021);
   U5374 : AO4 port map( A => n4474, B => n4349, C => n4710, D => n4631, Z => 
                           n4027);
   U5375 : AO4 port map( A => n4475, B => n4349, C => n4710, D => n4632, Z => 
                           n4034);
   U5376 : AO4 port map( A => n4476, B => n4349, C => n4710, D => n4633, Z => 
                           n4040);
   U5377 : AO4 port map( A => n4477, B => n4349, C => n4710, D => n4634, Z => 
                           n4046);
   U5378 : AO4 port map( A => n4478, B => n4349, C => n4710, D => n4635, Z => 
                           n4052);
   U5379 : AO4 port map( A => n4479, B => n4349, C => n4710, D => n4636, Z => 
                           n4058);
   U5380 : AO4 port map( A => n4480, B => n4349, C => n4710, D => n4637, Z => 
                           n4064);
   U5381 : AO4 port map( A => n4481, B => n4349, C => n4710, D => n4638, Z => 
                           n4070);
   U5382 : AO4 port map( A => n4482, B => n4349, C => n4710, D => n4639, Z => 
                           n4077);
   U5383 : AO4 port map( A => n4483, B => n4349, C => n4710, D => n4640, Z => 
                           n4083);
   U5384 : AO4 port map( A => n4484, B => n4349, C => n4710, D => n4641, Z => 
                           n4089);
   U5385 : AO4 port map( A => n4485, B => n4349, C => n4710, D => n4642, Z => 
                           n4095);
   U5386 : AO4 port map( A => n4486, B => n4349, C => n4710, D => n4643, Z => 
                           n4101);
   U5387 : AO4 port map( A => n4487, B => n4349, C => n4710, D => n4644, Z => 
                           n4108);
   U5388 : AO4 port map( A => n4488, B => n4349, C => n4710, D => n4645, Z => 
                           n4114);
   U5389 : AO4 port map( A => n4489, B => n4349, C => n4710, D => n4646, Z => 
                           n4120);
   U5390 : AO4 port map( A => n4490, B => n4349, C => n4710, D => n4647, Z => 
                           n4126);
   U5391 : AO4 port map( A => n4491, B => n4349, C => n4710, D => n4648, Z => 
                           n4133);
   U5392 : AO4 port map( A => n4492, B => n4349, C => n4710, D => n4649, Z => 
                           n4139);
   U5393 : AO4 port map( A => n4493, B => n4349, C => n4710, D => n4650, Z => 
                           n4145);
   U5394 : AO4 port map( A => n4494, B => n4349, C => n4710, D => n4651, Z => 
                           n4151);
   U5395 : AO4 port map( A => n4495, B => n4349, C => n4710, D => n4652, Z => 
                           n4158);
   U5396 : AO3 port map( A => n4462, B => n1467, C => n4843, D => n4349, Z => 
                           n1486);
   U5397 : AO7 port map( A => n4864, B => n4601, C => n1498, Z => n1491);
   U5398 : AO7 port map( A => n4713, B => n1398, C => n4850, Z => n1487);
   U5399 : ND3 port map( A => n4850, B => n4380, C => n1493, Z => n1489);
   U5400 : AO3 port map( A => n4350, B => n4377, C => n1491, D => n1492, Z => 
                           n1490);
   U5401 : ND3 port map( A => n4850, B => n4602, C => n1493, Z => n1494);
   U5402 : ND4 port map( A => n4855, B => n1491, C => n4579, D => n4384, Z => 
                           n1495);
   U5403 : IVDA port map( A => n1427, Y => n4584, Z => n4677);
   U5404 : IVDA port map( A => n1408, Y => n4585, Z => n4693);
   U5405 : NR4 port map( A => v_CALCULATION_CNTR_4_port, B => 
                           v_CALCULATION_CNTR_5_port, C => 
                           v_CALCULATION_CNTR_6_port, D => 
                           v_CALCULATION_CNTR_7_port, Z => n1499);
   U5406 : AO7 port map( A => n1386, B => n4713, C => n4850, Z => n105);
   U5407 : AO6 port map( A => n3955, B => n1387, C => n1353, Z => n1386);
   U5408 : AO3 port map( A => n4354, B => n4477, C => n293, D => n294, Z => 
                           n4050);
   U5409 : AO2 port map( A => n4496, B => n317, C => n318, D => n4382, Z => 
                           n293);
   U5410 : AO6 port map( A => n295, B => n4844, C => n296, Z => n294);
   U5411 : AO3 port map( A => n4354, B => n4478, C => n756, D => n757, Z => 
                           n4056);
   U5412 : AO2 port map( A => n4496, B => n783, C => n784, D => n4382, Z => 
                           n756);
   U5413 : AO6 port map( A => n758, B => n4844, C => n759, Z => n757);
   U5414 : AO3 port map( A => n4354, B => n4479, C => n1104, D => n1105, Z => 
                           n4062);
   U5415 : AO2 port map( A => n4496, B => n1148, C => n1149, D => n4382, Z => 
                           n1104);
   U5416 : AO6 port map( A => n1106, B => n4844, C => n1107, Z => n1105);
   U5417 : AO3 port map( A => n4354, B => n4480, C => n499, D => n500, Z => 
                           n4068);
   U5418 : AO2 port map( A => n4496, B => n517, C => n518, D => n4382, Z => 
                           n499);
   U5419 : AO6 port map( A => n501, B => n4844, C => n502, Z => n500);
   U5420 : AO4 port map( A => n978, B => n4711, C => n164, D => n979, Z => n969
                           );
   U5421 : AO4 port map( A => n162, B => n4711, C => n164, D => n165, Z => n149
                           );
   U5422 : AO3 port map( A => n4354, B => n4467, C => n930, D => n931, Z => 
                           n3989);
   U5423 : AO2 port map( A => n4496, B => n955, C => n956, D => n4382, Z => 
                           n930);
   U5424 : AO6 port map( A => n932, B => n4844, C => n933, Z => n931);
   U5425 : AO3 port map( A => n4354, B => n4468, C => n596, D => n597, Z => 
                           n3995);
   U5426 : AO2 port map( A => n4496, B => n614, C => n615, D => n4382, Z => 
                           n596);
   U5427 : AO6 port map( A => n598, B => n4844, C => n599, Z => n597);
   U5428 : AO3 port map( A => n4354, B => n4469, C => n326, D => n327, Z => 
                           n4001);
   U5429 : AO2 port map( A => n4496, B => n356, C => n357, D => n4382, Z => 
                           n326);
   U5430 : AO6 port map( A => n328, B => n4844, C => n329, Z => n327);
   U5431 : AO3 port map( A => n4354, B => n4470, C => n1164, D => n1165, Z => 
                           n4007);
   U5432 : AO2 port map( A => n4496, B => n1221, C => n1222, D => n4382, Z => 
                           n1164);
   U5433 : AO6 port map( A => n1166, B => n4844, C => n1167, Z => n1165);
   U5434 : AO3 port map( A => n4354, B => n4471, C => n835, D => n836, Z => 
                           n4013);
   U5435 : AO2 port map( A => n4496, B => n874, C => n875, D => n4382, Z => 
                           n835);
   U5436 : AO6 port map( A => n837, B => n4844, C => n838, Z => n836);
   U5437 : AO3 port map( A => n4354, B => n4472, C => n524, D => n525, Z => 
                           n4019);
   U5438 : AO2 port map( A => n4496, B => n552, C => n553, D => n4382, Z => 
                           n524);
   U5439 : AO6 port map( A => n526, B => n4844, C => n527, Z => n525);
   U5440 : AO3 port map( A => n4354, B => n4474, C => n563, D => n564, Z => 
                           n4031);
   U5441 : AO2 port map( A => n4496, B => n587, C => n588, D => n4382, Z => 
                           n563);
   U5442 : AO6 port map( A => n565, B => n4844, C => n566, Z => n564);
   U5443 : AO3 port map( A => n4354, B => n4475, C => n107, D => n108, Z => 
                           n4038);
   U5444 : AO2 port map( A => n4496, B => n135, C => n136, D => n4382, Z => 
                           n107);
   U5445 : AO6 port map( A => n109, B => n4844, C => n111, Z => n108);
   U5446 : AO3 port map( A => n4354, B => n4476, C => n793, D => n794, Z => 
                           n4044);
   U5447 : AO2 port map( A => n4496, B => n823, C => n824, D => n4382, Z => 
                           n793);
   U5448 : AO6 port map( A => n795, B => n4844, C => n796, Z => n794);
   U5449 : AO3 port map( A => n4354, B => n4481, C => n888, D => n889, Z => 
                           n4074);
   U5450 : AO2 port map( A => n4496, B => n918, C => n919, D => n4382, Z => 
                           n888);
   U5451 : AO6 port map( A => n890, B => n4844, C => n891, Z => n889);
   U5452 : AO3 port map( A => n4354, B => n4482, C => n425, D => n426, Z => 
                           n4081);
   U5453 : AO2 port map( A => n4496, B => n455, C => n456, D => n4382, Z => 
                           n425);
   U5454 : AO6 port map( A => n427, B => n4844, C => n428, Z => n426);
   U5455 : AO3 port map( A => n4354, B => n4483, C => n260, D => n261, Z => 
                           n4087);
   U5456 : AO2 port map( A => n4496, B => n284, C => n285, D => n4382, Z => 
                           n260);
   U5457 : AO6 port map( A => n262, B => n4844, C => n263, Z => n261);
   U5458 : AO3 port map( A => n4354, B => n4484, C => n466, D => n467, Z => 
                           n4093);
   U5459 : AO2 port map( A => n4496, B => n490, C => n491, D => n4382, Z => 
                           n466);
   U5460 : AO6 port map( A => n468, B => n4844, C => n469, Z => n467);
   U5461 : AO3 port map( A => n4354, B => n4485, C => n1065, D => n1066, Z => 
                           n4099);
   U5462 : AO2 port map( A => n4496, B => n1093, C => n1094, D => n4382, Z => 
                           n1065);
   U5463 : AO6 port map( A => n1067, B => n4844, C => n1068, Z => n1066);
   U5464 : AO3 port map( A => n4354, B => n4486, C => n731, D => n732, Z => 
                           n4105);
   U5465 : AO2 port map( A => n4496, B => n749, C => n750, D => n4382, Z => 
                           n731);
   U5466 : AO6 port map( A => n733, B => n4844, C => n734, Z => n732);
   U5467 : AO3 port map( A => n4354, B => n4487, C => n235, D => n236, Z => 
                           n4112);
   U5468 : AO2 port map( A => n4496, B => n253, C => n254, D => n4382, Z => 
                           n235);
   U5469 : AO6 port map( A => n237, B => n4844, C => n238, Z => n236);
   U5470 : AO3 port map( A => n4354, B => n4488, C => n1036, D => n1037, Z => 
                           n4118);
   U5471 : AO2 port map( A => n4496, B => n1057, C => n1058, D => n4382, Z => 
                           n1036);
   U5472 : AO6 port map( A => n1038, B => n4844, C => n1039, Z => n1037);
   U5473 : AO3 port map( A => n4354, B => n4489, C => n702, D => n703, Z => 
                           n4124);
   U5474 : AO2 port map( A => n4496, B => n723, C => n724, D => n4382, Z => 
                           n702);
   U5475 : AO6 port map( A => n704, B => n4844, C => n705, Z => n703);
   U5476 : AO3 port map( A => n4354, B => n4490, C => n392, D => n393, Z => 
                           n4130);
   U5477 : AO2 port map( A => n4496, B => n416, C => n417, D => n4382, Z => 
                           n392);
   U5478 : AO6 port map( A => n394, B => n4844, C => n395, Z => n393);
   U5479 : AO3 port map( A => n4354, B => n4491, C => n206, D => n207, Z => 
                           n4137);
   U5480 : AO2 port map( A => n4496, B => n227, C => n228, D => n4382, Z => 
                           n206);
   U5481 : AO6 port map( A => n208, B => n4844, C => n209, Z => n207);
   U5482 : AO3 port map( A => n4354, B => n4492, C => n1007, D => n1008, Z => 
                           n4143);
   U5483 : AO2 port map( A => n4496, B => n1027, C => n1028, D => n4382, Z => 
                           n1007);
   U5484 : AO6 port map( A => n1009, B => n4844, C => n1010, Z => n1008);
   U5485 : AO3 port map( A => n4354, B => n4493, C => n664, D => n665, Z => 
                           n4149);
   U5486 : AO2 port map( A => n4496, B => n692, C => n693, D => n4382, Z => 
                           n664);
   U5487 : AO6 port map( A => n666, B => n4844, C => n667, Z => n665);
   U5488 : AO3 port map( A => n4354, B => n4494, C => n367, D => n368, Z => 
                           n4155);
   U5489 : AO2 port map( A => n4496, B => n385, C => n386, D => n4382, Z => 
                           n367);
   U5490 : AO6 port map( A => n369, B => n4844, C => n370, Z => n368);
   U5491 : AO3 port map( A => n4354, B => n4495, C => n621, D => n622, Z => 
                           n4162);
   U5492 : AO2 port map( A => n4496, B => n652, C => n653, D => n4382, Z => 
                           n621);
   U5493 : AO6 port map( A => n623, B => n4844, C => n624, Z => n622);
   U5494 : AO4 port map( A => n1339, B => n4711, C => n164, D => n1340, Z => 
                           n1322);
   U5495 : AO3 port map( A => n4354, B => n4473, C => n1240, D => n1241, Z => 
                           n4025);
   U5496 : AO2 port map( A => n4496, B => n1297, C => n1298, D => n4382, Z => 
                           n1240);
   U5497 : AO6 port map( A => n1242, B => n4844, C => n1243, Z => n1241);
   U5498 : NR3 port map( A => n4860, B => RESET_I, C => n1353, Z => n1350);
   U5499 : AO7 port map( A => n3824, B => n1995, C => n1999, Z => n4171);
   U5500 : EO1 port map( A => n4389, B => n4786, C => n1991, D => n4903, Z => 
                           n1999);
   U5501 : AO7 port map( A => n3825, B => n1995, C => n4784, Z => n4172);
   U5502 : AO4 port map( A => n1991, B => n1651, C => n4706, D => n696, Z => 
                           n1997);
   U5503 : NR3 port map( A => n3951, B => n4845, C => n4852, Z => n1471);
   U5504 : AO4 port map( A => n3955, B => n4672, C => n4441, D => n1485, Z => 
                           n1459);
   U5505 : AO7 port map( A => n3954, B => n1459, C => CE_I, Z => n1482);
   U5506 : AO3 port map( A => n1621, B => n1917, C => n1931, D => n1932, Z => 
                           n4156);
   U5507 : AO3 port map( A => n4870, B => n1917, C => n1927, D => n1928, Z => 
                           n4163);
   U5508 : AO3 port map( A => n1603, B => n1917, C => n1918, D => n1919, Z => 
                           n4165);
   U5509 : AO7 port map( A => n3840, B => n2426, C => n2430, Z => n4187);
   U5510 : EO1 port map( A => n4389, B => n4757, C => n2422, D => n4911, Z => 
                           n2430);
   U5511 : AO7 port map( A => n3953, B => n1469, C => n1470, Z => n4286);
   U5512 : AO6 port map( A => n3952, B => n1474, C => n1475, Z => n1469);
   U5513 : ND4 port map( A => n3953, B => n1471, C => n4619, D => n4463, Z => 
                           n1470);
   U5514 : EON1 port map( A => n3950, B => n1477, C => n1471, D => n3950, Z => 
                           n4288);
   U5515 : NR4 port map( A => n4407, B => v_CALCULATION_CNTR_3_port, C => n4502
                           , D => n3809, Z => n3803);
   U5516 : ND2I port map( A => v_RAM_OUT0_19_port, B => n4501, Z => n2987);
   U5517 : ND2I port map( A => v_RAM_OUT0_3_port, B => n4500, Z => n3388);
   U5518 : AO3 port map( A => n4378, B => n2245, C => n2322, D => n2323, Z => 
                           n2321);
   U5519 : AO2 port map( A => n2032, B => n4702, C => n4701, D => n2133, Z => 
                           n2322);
   U5520 : AO3 port map( A => n1661, B => n2893, C => n3100, D => n3101, Z => 
                           n4202);
   U5521 : AO3 port map( A => n1651, B => n2893, C => n2971, D => n2972, Z => 
                           n4204);
   U5522 : AO3 port map( A => n1593, B => n1755, C => n1776, D => n1777, Z => 
                           n4247);
   U5523 : AO3 port map( A => n4911, B => n1755, C => n1763, D => n1764, Z => 
                           n4251);
   U5524 : AO3 port map( A => n1603, B => n1783, C => n1784, D => n1785, Z => 
                           n4261);
   U5525 : AO3 port map( A => n1651, B => n1811, C => n1816, D => n1817, Z => 
                           n4268);
   U5526 : ND2I port map( A => v_RAM_OUT0_27_port, B => n4508, Z => n2584);
   U5527 : AO4 port map( A => v_RAM_OUT0_12_port, B => n2234, C => n2402, D => 
                           n4404, Z => n1902);
   U5528 : AO4 port map( A => n3899, B => n4675, C => n3907, D => n4676, Z => 
                           n3795);
   U5529 : AO7 port map( A => n3811, B => n4672, C => n3799, Z => n3794);
   U5530 : AO2 port map( A => n1516, B => n4520, C => n1515, D => n4419, Z => 
                           n3799);
   U5531 : AO4 port map( A => n3900, B => n4675, C => n3908, D => n4676, Z => 
                           n3784);
   U5532 : AO7 port map( A => n3812, B => n4672, C => n3785, Z => n3783);
   U5533 : AO2 port map( A => n1516, B => n4570, C => n1515, D => n4445, Z => 
                           n3785);
   U5534 : AO4 port map( A => n3901, B => n4675, C => n3909, D => n4676, Z => 
                           n3773);
   U5535 : AO7 port map( A => n3813, B => n4672, C => n3774, Z => n3772);
   U5536 : AO2 port map( A => n1516, B => n4551, C => n1515, D => n4432, Z => 
                           n3774);
   U5537 : AO4 port map( A => n3902, B => n4675, C => n3910, D => n4676, Z => 
                           n3762);
   U5538 : AO7 port map( A => n3814, B => n4672, C => n3763, Z => n3761);
   U5539 : AO2 port map( A => n1516, B => n4552, C => n1515, D => n4455, Z => 
                           n3763);
   U5540 : AO4 port map( A => n3903, B => n4675, C => n3911, D => n4676, Z => 
                           n3751);
   U5541 : AO7 port map( A => n3815, B => n4672, C => n3752, Z => n3750);
   U5542 : AO2 port map( A => n1516, B => n4582, C => n1515, D => n4446, Z => 
                           n3752);
   U5543 : AO4 port map( A => n3904, B => n4675, C => n3912, D => n4676, Z => 
                           n3740);
   U5544 : AO7 port map( A => n3816, B => n4672, C => n3741, Z => n3739);
   U5545 : AO2 port map( A => n1516, B => n4415, C => n1515, D => n4580, Z => 
                           n3741);
   U5546 : AO4 port map( A => n3905, B => n4675, C => n3913, D => n4676, Z => 
                           n3729);
   U5547 : AO7 port map( A => n3817, B => n4672, C => n3730, Z => n3728);
   U5548 : AO2 port map( A => n1516, B => n4583, C => n1515, D => n4433, Z => 
                           n3730);
   U5549 : AO4 port map( A => n3906, B => n4675, C => n3914, D => n4676, Z => 
                           n3717);
   U5550 : AO7 port map( A => n3818, B => n4672, C => n3718, Z => n3716);
   U5551 : AO2 port map( A => n1516, B => n4420, C => n1515, D => n4581, Z => 
                           n3718);
   U5552 : AO2 port map( A => n5041, B => n2277, C => n4993, D => n5040, Z => 
                           n2274);
   U5553 : AO3 port map( A => n1621, B => n1783, C => n1795, D => n1796, Z => 
                           n4258);
   U5554 : AO3 port map( A => n1661, B => n1811, C => n1823, D => n1824, Z => 
                           n4266);
   U5555 : AO4 port map( A => n3951, B => n1480, C => n4845, D => n1481, Z => 
                           n4289);
   U5556 : AO3 port map( A => n3915, B => n4706, C => n3787, D => n3788, Z => 
                           n3958);
   U5557 : AO2 port map( A => n4709, B => n4519, C => n4673, D => DATA_O_0_port
                           , Z => n3788);
   U5558 : AO2 port map( A => n4366, B => n3789, C => n4708, D => n4545, Z => 
                           n3787);
   U5559 : ND4 port map( A => n3790, B => n3791, C => n3792, D => n3793, Z => 
                           n3789);
   U5560 : AO3 port map( A => n3916, B => n4706, C => n3776, D => n3777, Z => 
                           n3959);
   U5561 : AO2 port map( A => n4709, B => n4605, C => n4673, D => DATA_O_1_port
                           , Z => n3777);
   U5562 : AO2 port map( A => n4366, B => n3778, C => n4708, D => n4603, Z => 
                           n3776);
   U5563 : ND4 port map( A => n3779, B => n3780, C => n3781, D => n3782, Z => 
                           n3778);
   U5564 : AO3 port map( A => n3917, B => n4706, C => n3765, D => n3766, Z => 
                           n3960);
   U5565 : AO2 port map( A => n4709, B => n4532, C => n4673, D => DATA_O_2_port
                           , Z => n3766);
   U5566 : AO2 port map( A => n4366, B => n3767, C => n4708, D => n4517, Z => 
                           n3765);
   U5567 : ND4 port map( A => n3768, B => n3769, C => n3770, D => n3771, Z => 
                           n3767);
   U5568 : AO3 port map( A => n3918, B => n4706, C => n3754, D => n3755, Z => 
                           n3961);
   U5569 : AO2 port map( A => n4709, B => n4444, C => n4673, D => DATA_O_3_port
                           , Z => n3755);
   U5570 : AO2 port map( A => n4366, B => n3756, C => n4708, D => n4546, Z => 
                           n3754);
   U5571 : ND4 port map( A => n3757, B => n3758, C => n3759, D => n3760, Z => 
                           n3756);
   U5572 : AO3 port map( A => n3919, B => n4706, C => n3743, D => n3744, Z => 
                           n3962);
   U5573 : AO2 port map( A => n4709, B => n4550, C => n4673, D => DATA_O_4_port
                           , Z => n3744);
   U5574 : AO2 port map( A => n4366, B => n3745, C => n4708, D => n4547, Z => 
                           n3743);
   U5575 : ND4 port map( A => n3746, B => n3747, C => n3748, D => n3749, Z => 
                           n3745);
   U5576 : AO3 port map( A => n3920, B => n4706, C => n3732, D => n3733, Z => 
                           n3963);
   U5577 : AO2 port map( A => n4709, B => n4606, C => n4673, D => DATA_O_5_port
                           , Z => n3733);
   U5578 : AO2 port map( A => n4366, B => n3734, C => n4708, D => n4604, Z => 
                           n3732);
   U5579 : ND4 port map( A => n3735, B => n3736, C => n3737, D => n3738, Z => 
                           n3734);
   U5580 : AO3 port map( A => n3921, B => n4706, C => n3721, D => n3722, Z => 
                           n3964);
   U5581 : AO2 port map( A => n4709, B => n4431, C => n4673, D => DATA_O_6_port
                           , Z => n3722);
   U5582 : AO2 port map( A => n4366, B => n3723, C => n4708, D => n4416, Z => 
                           n3721);
   U5583 : ND4 port map( A => n3724, B => n3725, C => n3726, D => n3727, Z => 
                           n3723);
   U5584 : AO3 port map( A => n3922, B => n4706, C => n3705, D => n3706, Z => 
                           n3965);
   U5585 : AO2 port map( A => n4709, B => n4607, C => n4673, D => DATA_O_7_port
                           , Z => n3706);
   U5586 : AO2 port map( A => n4366, B => n3710, C => n4708, D => n4417, Z => 
                           n3705);
   U5587 : ND4 port map( A => n3712, B => n3713, C => n3714, D => n3715, Z => 
                           n3710);
   U5588 : AO2 port map( A => n4849, B => v_CALCULATION_CNTR_7_port, C => N2089
                           , D => n1450, Z => n1448);
   U5589 : AO2 port map( A => n4849, B => v_CALCULATION_CNTR_6_port, C => N2088
                           , D => n1450, Z => n1451);
   U5590 : AO2 port map( A => n4849, B => v_CALCULATION_CNTR_5_port, C => N2087
                           , D => n1450, Z => n1452);
   U5591 : NR4 port map( A => n2392, B => n4502, C => n3805, D => 
                           v_CALCULATION_CNTR_5_port, Z => n3802);
   U5592 : ND2I port map( A => v_RAM_OUT0_22_port, B => n4393, Z => n3019);
   U5593 : ND2I port map( A => v_RAM_OUT0_6_port, B => n4392, Z => n3420);
   U5594 : AO2 port map( A => v_RAM_OUT0_12_port, B => n4977, C => n4404, D => 
                           n2166, Z => n1876);
   U5595 : EON1 port map( A => v_RAM_OUT0_12_port, B => n2064, C => n4378, D =>
                           n2192, Z => n2265);
   U5596 : AO6 port map( A => n4674, B => n4530, C => n3801, Z => n3792);
   U5597 : AO4 port map( A => n3835, B => n1511, C => n3851, D => n1510, Z => 
                           n3801);
   U5598 : AO6 port map( A => n4674, B => n4548, C => n3786, Z => n3781);
   U5599 : AO4 port map( A => n3836, B => n1511, C => n3852, D => n1510, Z => 
                           n3786);
   U5600 : AO6 port map( A => n4674, B => n4549, C => n3775, Z => n3770);
   U5601 : AO4 port map( A => n3837, B => n1511, C => n3853, D => n1510, Z => 
                           n3775);
   U5602 : AO6 port map( A => n4674, B => n4531, C => n3764, Z => n3759);
   U5603 : AO4 port map( A => n3838, B => n1511, C => n3854, D => n1510, Z => 
                           n3764);
   U5604 : AO6 port map( A => n4674, B => n4594, C => n3753, Z => n3748);
   U5605 : AO4 port map( A => n3839, B => n1511, C => n3855, D => n1510, Z => 
                           n3753);
   U5606 : AO6 port map( A => n4674, B => n4514, C => n3742, Z => n3737);
   U5607 : AO4 port map( A => n3840, B => n1511, C => n3856, D => n1510, Z => 
                           n3742);
   U5608 : AO6 port map( A => n4674, B => n4526, C => n3731, Z => n3726);
   U5609 : AO4 port map( A => n3841, B => n1511, C => n3857, D => n1510, Z => 
                           n3731);
   U5610 : AO6 port map( A => n4674, B => n4518, C => n3719, Z => n3714);
   U5611 : AO4 port map( A => n3842, B => n1511, C => n3858, D => n1510, Z => 
                           n3719);
   U5612 : AO3 port map( A => n4359, B => n2245, C => n4906, D => n2259, Z => 
                           n2248);
   U5613 : AO6 port map( A => n4956, B => n4360, C => n2260, Z => n2259);
   U5614 : AO4 port map( A => n4361, B => n2261, C => n2262, D => n4707, Z => 
                           n2260);
   U5615 : AO6 port map( A => v_RAM_OUT0_11_port, B => n4391, C => n4966, Z => 
                           n2262);
   U5616 : AO4 port map( A => n3810, B => n4352, C => n3955, D => n1501, Z => 
                           n3957);
   U5617 : NR4 port map( A => n1516, B => n1517, C => n4564, D => n4452, Z => 
                           n1502);
   U5618 : NR4 port map( A => n1351, B => n1391, C => n4565, D => n1515, Z => 
                           n1503);
   U5619 : EON1 port map( A => n4502, B => n1454, C => N2086, D => n1450, Z => 
                           n4306);
   U5620 : EON1 port map( A => n4579, B => n1454, C => N2084, D => n1450, Z => 
                           n4308);
   U5621 : EOI port map( A => v_CALCULATION_CNTR_1_port, B => 
                           v_CALCULATION_CNTR_0_port, Z => N2083);
   U5622 : ND2I port map( A => v_RAM_OUT0_30_port, B => n4394, Z => n2617);
   U5623 : AO7 port map( A => n1474, B => n4849, C => n4441, Z => n3700);
   U5624 : ND4 port map( A => n3950, B => n4859, C => n4853, D => n3703, Z => 
                           n3701);
   U5625 : NR3 port map( A => n3953, B => n3952, C => n4713, Z => n3703);
   U5626 : EON1 port map( A => n4464, B => n4375, C => n4375, D => 
                           t_STATE_RAM0_1_0_port, Z => n3969);
   U5627 : EON1 port map( A => n4465, B => n4375, C => n4375, D => 
                           t_STATE_RAM0_1_16_port, Z => n3975);
   U5628 : EON1 port map( A => n4466, B => n4375, C => n4375, D => 
                           t_STATE_RAM0_1_8_port, Z => n3981);
   U5629 : EON1 port map( A => n4467, B => n4375, C => n4375, D => 
                           t_STATE_RAM0_1_17_port, Z => n3987);
   U5630 : EON1 port map( A => n4468, B => n4375, C => n4375, D => 
                           t_STATE_RAM0_1_25_port, Z => n3993);
   U5631 : EON1 port map( A => n4469, B => n4375, C => n4375, D => 
                           t_STATE_RAM0_1_3_port, Z => n3999);
   U5632 : EON1 port map( A => n4470, B => n4375, C => n4375, D => 
                           t_STATE_RAM0_1_11_port, Z => n4005);
   U5633 : EON1 port map( A => n4471, B => n4375, C => n4375, D => 
                           t_STATE_RAM0_1_19_port, Z => n4011);
   U5634 : EON1 port map( A => n4472, B => n4375, C => n4375, D => 
                           t_STATE_RAM0_1_27_port, Z => n4017);
   U5635 : EON1 port map( A => n4473, B => n4375, C => n4375, D => 
                           t_STATE_RAM0_1_10_port, Z => n4023);
   U5636 : EON1 port map( A => n4474, B => n4375, C => n4375, D => 
                           t_STATE_RAM0_1_26_port, Z => n4029);
   U5637 : EON1 port map( A => n4475, B => n4375, C => n4375, D => 
                           t_STATE_RAM0_1_9_port, Z => n4036);
   U5638 : EON1 port map( A => n4476, B => n4375, C => n4375, D => 
                           t_STATE_RAM0_1_1_port, Z => n4042);
   U5639 : EON1 port map( A => n4477, B => n4375, C => n4375, D => 
                           t_STATE_RAM0_1_4_port, Z => n4048);
   U5640 : EON1 port map( A => n4478, B => n4375, C => n4375, D => 
                           t_STATE_RAM0_1_20_port, Z => n4054);
   U5641 : EON1 port map( A => n4479, B => n4375, C => n4375, D => 
                           t_STATE_RAM0_1_12_port, Z => n4060);
   U5642 : EON1 port map( A => n4480, B => n4375, C => n4375, D => 
                           t_STATE_RAM0_1_28_port, Z => n4066);
   U5643 : EON1 port map( A => n4481, B => n4375, C => n4375, D => 
                           t_STATE_RAM0_1_18_port, Z => n4072);
   U5644 : EON1 port map( A => n4482, B => n4375, C => n4375, D => 
                           t_STATE_RAM0_1_2_port, Z => n4079);
   U5645 : EON1 port map( A => n4483, B => n4375, C => n4375, D => 
                           t_STATE_RAM0_1_5_port, Z => n4085);
   U5646 : EON1 port map( A => n4484, B => n4375, C => n4375, D => 
                           t_STATE_RAM0_1_29_port, Z => n4091);
   U5647 : EON1 port map( A => n4485, B => n4375, C => n4375, D => 
                           t_STATE_RAM0_1_13_port, Z => n4097);
   U5648 : EON1 port map( A => n4486, B => n4375, C => n4375, D => 
                           t_STATE_RAM0_1_21_port, Z => n4103);
   U5649 : EON1 port map( A => n4487, B => n4375, C => n4375, D => 
                           t_STATE_RAM0_1_6_port, Z => n4110);
   U5650 : EON1 port map( A => n4488, B => n4375, C => n4375, D => 
                           t_STATE_RAM0_1_14_port, Z => n4116);
   U5651 : EON1 port map( A => n4489, B => n4375, C => n4375, D => 
                           t_STATE_RAM0_1_22_port, Z => n4122);
   U5652 : EON1 port map( A => n4490, B => n4375, C => n4375, D => 
                           t_STATE_RAM0_1_30_port, Z => n4128);
   U5653 : EON1 port map( A => n4491, B => n4375, C => n4375, D => 
                           t_STATE_RAM0_1_7_port, Z => n4135);
   U5654 : EON1 port map( A => n4492, B => n4375, C => n4375, D => 
                           t_STATE_RAM0_1_15_port, Z => n4141);
   U5655 : EON1 port map( A => n4493, B => n4375, C => n4375, D => 
                           t_STATE_RAM0_1_23_port, Z => n4147);
   U5656 : EON1 port map( A => n4494, B => n4375, C => n4375, D => 
                           t_STATE_RAM0_1_31_port, Z => n4153);
   U5657 : EON1 port map( A => n4495, B => n4375, C => n4375, D => 
                           t_STATE_RAM0_1_24_port, Z => n4160);
   U5658 : AO3 port map( A => n3954, B => n1454, C => n3806, D => n3807, Z => 
                           n4290);
   U5659 : ND4 port map( A => CE_I, B => n4850, C => n4840, D => n4527, Z => 
                           n3807);
   U5660 : AO7 port map( A => n3955, B => n4672, C => n1474, Z => n3806);
   U5661 : AO3 port map( A => n1392, B => n3944, C => n1393, D => n1394, Z => 
                           n4298);
   U5662 : AO7 port map( A => n4841, B => RESET_I, C => n1392, Z => n1393);
   U5663 : AO7 port map( A => n3949, B => n4713, C => n4843, Z => n1392);
   U5664 : EON1 port map( A => n4464, B => n4358, C => n4358, D => 
                           t_STATE_RAM0_2_0_port, Z => n3968);
   U5665 : EON1 port map( A => n4466, B => n4358, C => n4358, D => 
                           t_STATE_RAM0_2_8_port, Z => n3980);
   U5666 : EON1 port map( A => n4468, B => n4358, C => n4358, D => 
                           t_STATE_RAM0_2_25_port, Z => n3992);
   U5667 : EON1 port map( A => n4469, B => n4358, C => n4358, D => 
                           t_STATE_RAM0_2_3_port, Z => n3998);
   U5668 : EON1 port map( A => n4472, B => n4358, C => n4358, D => 
                           t_STATE_RAM0_2_27_port, Z => n4016);
   U5669 : EON1 port map( A => n4474, B => n4358, C => n4358, D => 
                           t_STATE_RAM0_2_26_port, Z => n4028);
   U5670 : EON1 port map( A => n4475, B => n4358, C => n4358, D => 
                           t_STATE_RAM0_2_9_port, Z => n4035);
   U5671 : EON1 port map( A => n4477, B => n4358, C => n4358, D => 
                           t_STATE_RAM0_2_4_port, Z => n4047);
   U5672 : EON1 port map( A => n4480, B => n4358, C => n4358, D => 
                           t_STATE_RAM0_2_28_port, Z => n4065);
   U5673 : EON1 port map( A => n4482, B => n4358, C => n4358, D => 
                           t_STATE_RAM0_2_2_port, Z => n4078);
   U5674 : EON1 port map( A => n4483, B => n4358, C => n4358, D => 
                           t_STATE_RAM0_2_5_port, Z => n4084);
   U5675 : EON1 port map( A => n4484, B => n4358, C => n4358, D => 
                           t_STATE_RAM0_2_29_port, Z => n4090);
   U5676 : EON1 port map( A => n4487, B => n4358, C => n4358, D => 
                           t_STATE_RAM0_2_6_port, Z => n4109);
   U5677 : EON1 port map( A => n4490, B => n4358, C => n4358, D => 
                           t_STATE_RAM0_2_30_port, Z => n4127);
   U5678 : EON1 port map( A => n4491, B => n4358, C => n4358, D => 
                           t_STATE_RAM0_2_7_port, Z => n4134);
   U5679 : EON1 port map( A => n4494, B => n4358, C => n4358, D => 
                           t_STATE_RAM0_2_31_port, Z => n4152);
   U5680 : AO3 port map( A => n1392, B => n3941, C => n1393, D => n1395, Z => 
                           n4293);
   U5681 : AO3 port map( A => n1392, B => n3942, C => n1393, D => n1396, Z => 
                           n4294);
   U5682 : AO7 port map( A => n1392, B => n3943, C => n1397, Z => n4295);
   U5683 : ND4 port map( A => N200, B => n1392, C => n1398, D => n4850, Z => 
                           n1397);
   U5684 : AO3 port map( A => n4653, B => n1392, C => n1393, D => n1399, Z => 
                           n4296);
   U5685 : AO3 port map( A => n4620, B => n1392, C => n1393, D => n1400, Z => 
                           n4297);
   U5686 : ND4 port map( A => CE_I, B => n1499, C => n4579, D => n4384, Z => 
                           n1493);
   U5687 : AO3 port map( A => n4381, B => n4621, C => n100, D => n101, Z => 
                           n3966);
   U5688 : AO2 port map( A => t_STATE_RAM0_0_0_port, B => n4351, C => 
                           t_STATE_RAM0_2_0_port, D => n4350, Z => n100);
   U5689 : AO2 port map( A => t_STATE_RAM0_1_0_port, B => n4377, C => 
                           v_RAM_OUT0_0_port, D => n4713, Z => n101);
   U5690 : EON1 port map( A => n4464, B => n4376, C => n4376, D => 
                           t_STATE_RAM0_0_0_port, Z => n3970);
   U5691 : AO3 port map( A => n4381, B => n4622, C => n79, D => n80, Z => n3972
                           );
   U5692 : AO2 port map( A => t_STATE_RAM0_0_16_port, B => n4351, C => 
                           t_STATE_RAM0_2_16_port, D => n4350, Z => n79);
   U5693 : AO2 port map( A => t_STATE_RAM0_1_16_port, B => n4377, C => 
                           v_RAM_OUT0_16_port, D => n4713, Z => n80);
   U5694 : EON1 port map( A => n4465, B => n4358, C => n4358, D => 
                           t_STATE_RAM0_2_16_port, Z => n3974);
   U5695 : EON1 port map( A => n4465, B => n4376, C => n4376, D => 
                           t_STATE_RAM0_0_16_port, Z => n3976);
   U5696 : AO3 port map( A => n4381, B => n4623, C => n10, D => n11, Z => n3978
                           );
   U5697 : AO2 port map( A => t_STATE_RAM0_0_8_port, B => n4351, C => 
                           t_STATE_RAM0_2_8_port, D => n4350, Z => n10);
   U5698 : AO2 port map( A => t_STATE_RAM0_1_8_port, B => n4377, C => 
                           v_RAM_OUT0_8_port, D => n4713, Z => n11);
   U5699 : EON1 port map( A => n4466, B => n4376, C => n4376, D => 
                           t_STATE_RAM0_0_8_port, Z => n3982);
   U5700 : AO3 port map( A => n4381, B => n4624, C => n76, D => n77, Z => n3984
                           );
   U5701 : AO2 port map( A => t_STATE_RAM0_0_17_port, B => n4351, C => 
                           t_STATE_RAM0_2_17_port, D => n4350, Z => n76);
   U5702 : AO2 port map( A => t_STATE_RAM0_1_17_port, B => n4377, C => 
                           v_RAM_OUT0_17_port, D => n4713, Z => n77);
   U5703 : EON1 port map( A => n4467, B => n4358, C => n4358, D => 
                           t_STATE_RAM0_2_17_port, Z => n3986);
   U5704 : EON1 port map( A => n4467, B => n4376, C => n4376, D => 
                           t_STATE_RAM0_0_17_port, Z => n3988);
   U5705 : AO3 port map( A => n4381, B => n4625, C => n49, D => n50, Z => n3990
                           );
   U5706 : AO2 port map( A => t_STATE_RAM0_0_25_port, B => n4351, C => 
                           t_STATE_RAM0_2_25_port, D => n4350, Z => n49);
   U5707 : AO2 port map( A => t_STATE_RAM0_1_25_port, B => n4377, C => 
                           v_RAM_OUT0_25_port, D => n4713, Z => n50);
   U5708 : EON1 port map( A => n4468, B => n4376, C => n4376, D => 
                           t_STATE_RAM0_0_25_port, Z => n3994);
   U5709 : AO3 port map( A => n4381, B => n4626, C => n25, D => n26, Z => n3996
                           );
   U5710 : AO2 port map( A => t_STATE_RAM0_0_3_port, B => n4351, C => 
                           t_STATE_RAM0_2_3_port, D => n4350, Z => n25);
   U5711 : AO2 port map( A => t_STATE_RAM0_1_3_port, B => n4377, C => 
                           v_RAM_OUT0_3_port, D => n4713, Z => n26);
   U5712 : EON1 port map( A => n4469, B => n4376, C => n4376, D => 
                           t_STATE_RAM0_0_3_port, Z => n4000);
   U5713 : AO3 port map( A => n4381, B => n4627, C => n94, D => n95, Z => n4002
                           );
   U5714 : AO2 port map( A => t_STATE_RAM0_0_11_port, B => n4351, C => 
                           t_STATE_RAM0_2_11_port, D => n4350, Z => n94);
   U5715 : AO2 port map( A => t_STATE_RAM0_1_11_port, B => n4377, C => 
                           v_RAM_OUT0_11_port, D => n4713, Z => n95);
   U5716 : EON1 port map( A => n4470, B => n4358, C => n4358, D => 
                           t_STATE_RAM0_2_11_port, Z => n4004);
   U5717 : EON1 port map( A => n4470, B => n4376, C => n4376, D => 
                           t_STATE_RAM0_0_11_port, Z => n4006);
   U5718 : AO3 port map( A => n4381, B => n4628, C => n70, D => n71, Z => n4008
                           );
   U5719 : AO2 port map( A => t_STATE_RAM0_0_19_port, B => n4351, C => 
                           t_STATE_RAM0_2_19_port, D => n4350, Z => n70);
   U5720 : AO2 port map( A => t_STATE_RAM0_1_19_port, B => n4377, C => 
                           v_RAM_OUT0_19_port, D => n4713, Z => n71);
   U5721 : EON1 port map( A => n4471, B => n4358, C => n4358, D => 
                           t_STATE_RAM0_2_19_port, Z => n4010);
   U5722 : EON1 port map( A => n4471, B => n4376, C => n4376, D => 
                           t_STATE_RAM0_0_19_port, Z => n4012);
   U5723 : AO3 port map( A => n4381, B => n4629, C => n43, D => n44, Z => n4014
                           );
   U5724 : AO2 port map( A => t_STATE_RAM0_0_27_port, B => n4351, C => 
                           t_STATE_RAM0_2_27_port, D => n4350, Z => n43);
   U5725 : AO2 port map( A => t_STATE_RAM0_1_27_port, B => n4377, C => 
                           v_RAM_OUT0_27_port, D => n4713, Z => n44);
   U5726 : EON1 port map( A => n4472, B => n4376, C => n4376, D => 
                           t_STATE_RAM0_0_27_port, Z => n4018);
   U5727 : AO3 port map( A => n4381, B => n4630, C => n97, D => n98, Z => n4020
                           );
   U5728 : AO2 port map( A => t_STATE_RAM0_0_10_port, B => n4351, C => 
                           t_STATE_RAM0_2_10_port, D => n4350, Z => n97);
   U5729 : AO2 port map( A => t_STATE_RAM0_1_10_port, B => n4377, C => 
                           v_RAM_OUT0_10_port, D => n4713, Z => n98);
   U5730 : EON1 port map( A => n4473, B => n4358, C => n4358, D => 
                           t_STATE_RAM0_2_10_port, Z => n4022);
   U5731 : EON1 port map( A => n4473, B => n4376, C => n4376, D => 
                           t_STATE_RAM0_0_10_port, Z => n4024);
   U5732 : AO3 port map( A => n4381, B => n4631, C => n46, D => n47, Z => n4026
                           );
   U5733 : AO2 port map( A => t_STATE_RAM0_0_26_port, B => n4351, C => 
                           t_STATE_RAM0_2_26_port, D => n4350, Z => n46);
   U5734 : AO2 port map( A => t_STATE_RAM0_1_26_port, B => n4377, C => 
                           v_RAM_OUT0_26_port, D => n4713, Z => n47);
   U5735 : EON1 port map( A => n4474, B => n4376, C => n4376, D => 
                           t_STATE_RAM0_0_26_port, Z => n4030);
   U5736 : AO3 port map( A => n4381, B => n4632, C => n3, D => n4, Z => n4033);
   U5737 : AO2 port map( A => t_STATE_RAM0_0_9_port, B => n4351, C => 
                           t_STATE_RAM0_2_9_port, D => n4350, Z => n3);
   U5738 : AO2 port map( A => t_STATE_RAM0_1_9_port, B => n4377, C => 
                           v_RAM_OUT0_9_port, D => n4713, Z => n4);
   U5739 : EON1 port map( A => n4475, B => n4376, C => n4376, D => 
                           t_STATE_RAM0_0_9_port, Z => n4037);
   U5740 : AO3 port map( A => n4381, B => n4633, C => n67, D => n68, Z => n4039
                           );
   U5741 : AO2 port map( A => t_STATE_RAM0_0_1_port, B => n4351, C => 
                           t_STATE_RAM0_2_1_port, D => n4350, Z => n67);
   U5742 : AO2 port map( A => t_STATE_RAM0_1_1_port, B => n4377, C => 
                           v_RAM_OUT0_1_port, D => n4713, Z => n68);
   U5743 : EON1 port map( A => n4476, B => n4358, C => n4358, D => 
                           t_STATE_RAM0_2_1_port, Z => n4041);
   U5744 : EON1 port map( A => n4476, B => n4376, C => n4376, D => 
                           t_STATE_RAM0_0_1_port, Z => n4043);
   U5745 : AO3 port map( A => n4381, B => n4634, C => n22, D => n23, Z => n4045
                           );
   U5746 : AO2 port map( A => t_STATE_RAM0_0_4_port, B => n4351, C => 
                           t_STATE_RAM0_2_4_port, D => n4350, Z => n22);
   U5747 : AO2 port map( A => t_STATE_RAM0_1_4_port, B => n4377, C => 
                           v_RAM_OUT0_4_port, D => n4713, Z => n23);
   U5748 : EON1 port map( A => n4477, B => n4376, C => n4376, D => 
                           t_STATE_RAM0_0_4_port, Z => n4049);
   U5749 : AO3 port map( A => n4381, B => n4635, C => n64, D => n65, Z => n4051
                           );
   U5750 : AO2 port map( A => t_STATE_RAM0_0_20_port, B => n4351, C => 
                           t_STATE_RAM0_2_20_port, D => n4350, Z => n64);
   U5751 : AO2 port map( A => t_STATE_RAM0_1_20_port, B => n4377, C => 
                           v_RAM_OUT0_20_port, D => n4713, Z => n65);
   U5752 : EON1 port map( A => n4478, B => n4358, C => n4358, D => 
                           t_STATE_RAM0_2_20_port, Z => n4053);
   U5753 : EON1 port map( A => n4478, B => n4376, C => n4376, D => 
                           t_STATE_RAM0_0_20_port, Z => n4055);
   U5754 : AO3 port map( A => n4381, B => n4636, C => n91, D => n92, Z => n4057
                           );
   U5755 : AO2 port map( A => t_STATE_RAM0_0_12_port, B => n4351, C => 
                           t_STATE_RAM0_2_12_port, D => n4350, Z => n91);
   U5756 : AO2 port map( A => t_STATE_RAM0_1_12_port, B => n4377, C => 
                           v_RAM_OUT0_12_port, D => n4713, Z => n92);
   U5757 : EON1 port map( A => n4479, B => n4358, C => n4358, D => 
                           t_STATE_RAM0_2_12_port, Z => n4059);
   U5758 : EON1 port map( A => n4479, B => n4376, C => n4376, D => 
                           t_STATE_RAM0_0_12_port, Z => n4061);
   U5759 : AO3 port map( A => n4381, B => n4637, C => n40, D => n41, Z => n4063
                           );
   U5760 : AO2 port map( A => t_STATE_RAM0_0_28_port, B => n4351, C => 
                           t_STATE_RAM0_2_28_port, D => n4350, Z => n40);
   U5761 : AO2 port map( A => t_STATE_RAM0_1_28_port, B => n4377, C => 
                           v_RAM_OUT0_28_port, D => n4713, Z => n41);
   U5762 : EON1 port map( A => n4480, B => n4376, C => n4376, D => 
                           t_STATE_RAM0_0_28_port, Z => n4067);
   U5763 : AO3 port map( A => n4381, B => n4638, C => n73, D => n74, Z => n4069
                           );
   U5764 : AO2 port map( A => t_STATE_RAM0_0_18_port, B => n4351, C => 
                           t_STATE_RAM0_2_18_port, D => n4350, Z => n73);
   U5765 : AO2 port map( A => t_STATE_RAM0_1_18_port, B => n4377, C => 
                           v_RAM_OUT0_18_port, D => n4713, Z => n74);
   U5766 : EON1 port map( A => n4481, B => n4358, C => n4358, D => 
                           t_STATE_RAM0_2_18_port, Z => n4071);
   U5767 : EON1 port map( A => n4481, B => n4376, C => n4376, D => 
                           t_STATE_RAM0_0_18_port, Z => n4073);
   U5768 : AO3 port map( A => n4381, B => n4639, C => n34, D => n35, Z => n4076
                           );
   U5769 : AO2 port map( A => t_STATE_RAM0_0_2_port, B => n4351, C => 
                           t_STATE_RAM0_2_2_port, D => n4350, Z => n34);
   U5770 : AO2 port map( A => t_STATE_RAM0_1_2_port, B => n4377, C => 
                           v_RAM_OUT0_2_port, D => n4713, Z => n35);
   U5771 : EON1 port map( A => n4482, B => n4376, C => n4376, D => 
                           t_STATE_RAM0_0_2_port, Z => n4080);
   U5772 : AO3 port map( A => n4381, B => n4640, C => n19, D => n20, Z => n4082
                           );
   U5773 : AO2 port map( A => t_STATE_RAM0_0_5_port, B => n4351, C => 
                           t_STATE_RAM0_2_5_port, D => n4350, Z => n19);
   U5774 : AO2 port map( A => t_STATE_RAM0_1_5_port, B => n4377, C => 
                           v_RAM_OUT0_5_port, D => n4713, Z => n20);
   U5775 : EON1 port map( A => n4483, B => n4376, C => n4376, D => 
                           t_STATE_RAM0_0_5_port, Z => n4086);
   U5776 : AO3 port map( A => n4381, B => n4641, C => n37, D => n38, Z => n4088
                           );
   U5777 : AO2 port map( A => t_STATE_RAM0_0_29_port, B => n4351, C => 
                           t_STATE_RAM0_2_29_port, D => n4350, Z => n37);
   U5778 : AO2 port map( A => t_STATE_RAM0_1_29_port, B => n4377, C => 
                           v_RAM_OUT0_29_port, D => n4713, Z => n38);
   U5779 : EON1 port map( A => n4484, B => n4376, C => n4376, D => 
                           t_STATE_RAM0_0_29_port, Z => n4092);
   U5780 : AO3 port map( A => n4381, B => n4642, C => n88, D => n89, Z => n4094
                           );
   U5781 : AO2 port map( A => t_STATE_RAM0_0_13_port, B => n4351, C => 
                           t_STATE_RAM0_2_13_port, D => n4350, Z => n88);
   U5782 : AO2 port map( A => t_STATE_RAM0_1_13_port, B => n4377, C => 
                           v_RAM_OUT0_13_port, D => n4713, Z => n89);
   U5783 : EON1 port map( A => n4485, B => n4358, C => n4358, D => 
                           t_STATE_RAM0_2_13_port, Z => n4096);
   U5784 : EON1 port map( A => n4485, B => n4376, C => n4376, D => 
                           t_STATE_RAM0_0_13_port, Z => n4098);
   U5785 : AO3 port map( A => n4381, B => n4643, C => n61, D => n62, Z => n4100
                           );
   U5786 : AO2 port map( A => t_STATE_RAM0_0_21_port, B => n4351, C => 
                           t_STATE_RAM0_2_21_port, D => n4350, Z => n61);
   U5787 : AO2 port map( A => t_STATE_RAM0_1_21_port, B => n4377, C => 
                           v_RAM_OUT0_21_port, D => n4713, Z => n62);
   U5788 : EON1 port map( A => n4486, B => n4358, C => n4358, D => 
                           t_STATE_RAM0_2_21_port, Z => n4102);
   U5789 : EON1 port map( A => n4486, B => n4376, C => n4376, D => 
                           t_STATE_RAM0_0_21_port, Z => n4104);
   U5790 : AO3 port map( A => n4381, B => n4644, C => n16, D => n17, Z => n4107
                           );
   U5791 : AO2 port map( A => t_STATE_RAM0_0_6_port, B => n4351, C => 
                           t_STATE_RAM0_2_6_port, D => n4350, Z => n16);
   U5792 : AO2 port map( A => t_STATE_RAM0_1_6_port, B => n4377, C => 
                           v_RAM_OUT0_6_port, D => n4713, Z => n17);
   U5793 : EON1 port map( A => n4487, B => n4376, C => n4376, D => 
                           t_STATE_RAM0_0_6_port, Z => n4111);
   U5794 : AO3 port map( A => n4381, B => n4645, C => n85, D => n86, Z => n4113
                           );
   U5795 : AO2 port map( A => t_STATE_RAM0_0_14_port, B => n4351, C => 
                           t_STATE_RAM0_2_14_port, D => n4350, Z => n85);
   U5796 : AO2 port map( A => t_STATE_RAM0_1_14_port, B => n4377, C => 
                           v_RAM_OUT0_14_port, D => n4713, Z => n86);
   U5797 : EON1 port map( A => n4488, B => n4358, C => n4358, D => 
                           t_STATE_RAM0_2_14_port, Z => n4115);
   U5798 : EON1 port map( A => n4488, B => n4376, C => n4376, D => 
                           t_STATE_RAM0_0_14_port, Z => n4117);
   U5799 : AO3 port map( A => n4381, B => n4646, C => n58, D => n59, Z => n4119
                           );
   U5800 : AO2 port map( A => t_STATE_RAM0_0_22_port, B => n4351, C => 
                           t_STATE_RAM0_2_22_port, D => n4350, Z => n58);
   U5801 : AO2 port map( A => t_STATE_RAM0_1_22_port, B => n4377, C => 
                           v_RAM_OUT0_22_port, D => n4713, Z => n59);
   U5802 : EON1 port map( A => n4489, B => n4358, C => n4358, D => 
                           t_STATE_RAM0_2_22_port, Z => n4121);
   U5803 : EON1 port map( A => n4489, B => n4376, C => n4376, D => 
                           t_STATE_RAM0_0_22_port, Z => n4123);
   U5804 : AO3 port map( A => n4381, B => n4647, C => n31, D => n32, Z => n4125
                           );
   U5805 : AO2 port map( A => t_STATE_RAM0_0_30_port, B => n4351, C => 
                           t_STATE_RAM0_2_30_port, D => n4350, Z => n31);
   U5806 : AO2 port map( A => t_STATE_RAM0_1_30_port, B => n4377, C => 
                           v_RAM_OUT0_30_port, D => n4713, Z => n32);
   U5807 : EON1 port map( A => n4490, B => n4376, C => n4376, D => 
                           t_STATE_RAM0_0_30_port, Z => n4129);
   U5808 : AO3 port map( A => n4381, B => n4648, C => n13, D => n14, Z => n4132
                           );
   U5809 : AO2 port map( A => t_STATE_RAM0_0_7_port, B => n4351, C => 
                           t_STATE_RAM0_2_7_port, D => n4350, Z => n13);
   U5810 : AO2 port map( A => t_STATE_RAM0_1_7_port, B => n4377, C => 
                           v_RAM_OUT0_7_port, D => n4713, Z => n14);
   U5811 : EON1 port map( A => n4491, B => n4376, C => n4376, D => 
                           t_STATE_RAM0_0_7_port, Z => n4136);
   U5812 : AO3 port map( A => n4381, B => n4649, C => n82, D => n83, Z => n4138
                           );
   U5813 : AO2 port map( A => t_STATE_RAM0_0_15_port, B => n4351, C => 
                           t_STATE_RAM0_2_15_port, D => n4350, Z => n82);
   U5814 : AO2 port map( A => t_STATE_RAM0_1_15_port, B => n4377, C => 
                           v_RAM_OUT0_15_port, D => n4713, Z => n83);
   U5815 : EON1 port map( A => n4492, B => n4358, C => n4358, D => 
                           t_STATE_RAM0_2_15_port, Z => n4140);
   U5816 : EON1 port map( A => n4492, B => n4376, C => n4376, D => 
                           t_STATE_RAM0_0_15_port, Z => n4142);
   U5817 : AO3 port map( A => n4381, B => n4650, C => n55, D => n56, Z => n4144
                           );
   U5818 : AO2 port map( A => t_STATE_RAM0_0_23_port, B => n4351, C => 
                           t_STATE_RAM0_2_23_port, D => n4350, Z => n55);
   U5819 : AO2 port map( A => t_STATE_RAM0_1_23_port, B => n4377, C => 
                           v_RAM_OUT0_23_port, D => n4713, Z => n56);
   U5820 : EON1 port map( A => n4493, B => n4358, C => n4358, D => 
                           t_STATE_RAM0_2_23_port, Z => n4146);
   U5821 : EON1 port map( A => n4493, B => n4376, C => n4376, D => 
                           t_STATE_RAM0_0_23_port, Z => n4148);
   U5822 : AO3 port map( A => n4381, B => n4651, C => n28, D => n29, Z => n4150
                           );
   U5823 : AO2 port map( A => t_STATE_RAM0_0_31_port, B => n4351, C => 
                           t_STATE_RAM0_2_31_port, D => n4350, Z => n28);
   U5824 : AO2 port map( A => t_STATE_RAM0_1_31_port, B => n4377, C => 
                           v_RAM_OUT0_31_port, D => n4713, Z => n29);
   U5825 : EON1 port map( A => n4494, B => n4376, C => n4376, D => 
                           t_STATE_RAM0_0_31_port, Z => n4154);
   U5826 : AO3 port map( A => n4381, B => n4652, C => n52, D => n53, Z => n4157
                           );
   U5827 : AO2 port map( A => t_STATE_RAM0_0_24_port, B => n4351, C => 
                           t_STATE_RAM0_2_24_port, D => n4350, Z => n52);
   U5828 : AO2 port map( A => t_STATE_RAM0_1_24_port, B => n4377, C => 
                           v_RAM_OUT0_24_port, D => n4713, Z => n53);
   U5829 : EON1 port map( A => n4495, B => n4358, C => n4358, D => 
                           t_STATE_RAM0_2_24_port, Z => n4159);
   U5830 : EON1 port map( A => n4495, B => n4376, C => n4376, D => 
                           t_STATE_RAM0_0_24_port, Z => n4161);
   U5831 : AO2 port map( A => n4677, B => v_DATA_COLUMN_23_port, C => DATA_I(7)
                           , D => n4584, Z => n1426);
   U5832 : AO2 port map( A => n4677, B => v_DATA_COLUMN_22_port, C => DATA_I(6)
                           , D => n4584, Z => n1429);
   U5833 : AO2 port map( A => n4677, B => v_DATA_COLUMN_21_port, C => DATA_I(5)
                           , D => n4584, Z => n1430);
   U5834 : AO2 port map( A => n4677, B => v_DATA_COLUMN_20_port, C => DATA_I(4)
                           , D => n4584, Z => n1431);
   U5835 : AO2 port map( A => n4677, B => v_DATA_COLUMN_19_port, C => DATA_I(3)
                           , D => n4584, Z => n1433);
   U5836 : AO2 port map( A => n4677, B => v_DATA_COLUMN_18_port, C => DATA_I(2)
                           , D => n4584, Z => n1434);
   U5837 : AO2 port map( A => n4677, B => v_DATA_COLUMN_17_port, C => DATA_I(1)
                           , D => n4584, Z => n1435);
   U5838 : AO2 port map( A => n4677, B => v_DATA_COLUMN_16_port, C => DATA_I(0)
                           , D => n4584, Z => n1436);
   U5839 : IVDA port map( A => n1404, Y => n4589, Z => n4692);
   U5840 : IVDA port map( A => n1415, Y => n4586, Z => n4694);
   U5841 : AO3 port map( A => CE_I, B => n4426, C => n1445, D => n4677, Z => 
                           n4337);
   U5842 : AO2 port map( A => n4693, B => v_DATA_COLUMN_7_port, C => n4585, D 
                           => DATA_I(7), Z => n1407);
   U5843 : AO2 port map( A => n4693, B => v_DATA_COLUMN_6_port, C => n4585, D 
                           => DATA_I(6), Z => n1410);
   U5844 : AO2 port map( A => n4693, B => v_DATA_COLUMN_5_port, C => n4585, D 
                           => DATA_I(5), Z => n1411);
   U5845 : AO2 port map( A => n4693, B => v_DATA_COLUMN_4_port, C => n4585, D 
                           => DATA_I(4), Z => n1412);
   U5846 : AO2 port map( A => n4693, B => v_DATA_COLUMN_3_port, C => n4585, D 
                           => DATA_I(3), Z => n1413);
   U5847 : AO2 port map( A => n4693, B => v_DATA_COLUMN_2_port, C => n4585, D 
                           => DATA_I(2), Z => n1418);
   U5848 : AO2 port map( A => n4693, B => v_DATA_COLUMN_1_port, C => DATA_I(1),
                           D => n4585, Z => n1432);
   U5849 : AO2 port map( A => n4693, B => v_DATA_COLUMN_0_port, C => DATA_I(0),
                           D => n4585, Z => n1443);
   U5850 : AO2 port map( A => n4692, B => v_DATA_COLUMN_15_port, C => n4589, D 
                           => DATA_I(7), Z => n1437);
   U5851 : AO2 port map( A => n4692, B => v_DATA_COLUMN_14_port, C => n4589, D 
                           => DATA_I(6), Z => n1438);
   U5852 : AO2 port map( A => n4692, B => v_DATA_COLUMN_13_port, C => n4589, D 
                           => DATA_I(5), Z => n1439);
   U5853 : AO2 port map( A => n4692, B => v_DATA_COLUMN_12_port, C => n4589, D 
                           => DATA_I(4), Z => n1440);
   U5854 : AO2 port map( A => n4692, B => v_DATA_COLUMN_11_port, C => n4589, D 
                           => DATA_I(3), Z => n1441);
   U5855 : AO2 port map( A => n4692, B => v_DATA_COLUMN_10_port, C => n4589, D 
                           => DATA_I(2), Z => n1442);
   U5856 : AO2 port map( A => n4692, B => v_DATA_COLUMN_9_port, C => n4589, D 
                           => DATA_I(1), Z => n1403);
   U5857 : AO2 port map( A => n4692, B => v_DATA_COLUMN_8_port, C => n4589, D 
                           => DATA_I(0), Z => n1406);
   U5858 : AO2 port map( A => n4694, B => v_DATA_COLUMN_31_port, C => DATA_I(7)
                           , D => n4586, Z => n1414);
   U5859 : AO2 port map( A => n4694, B => v_DATA_COLUMN_30_port, C => DATA_I(6)
                           , D => n4586, Z => n1417);
   U5860 : AO2 port map( A => n4694, B => v_DATA_COLUMN_29_port, C => DATA_I(5)
                           , D => n4586, Z => n1419);
   U5861 : AO2 port map( A => n4694, B => v_DATA_COLUMN_28_port, C => DATA_I(4)
                           , D => n4586, Z => n1420);
   U5862 : AO2 port map( A => n4694, B => v_DATA_COLUMN_27_port, C => DATA_I(3)
                           , D => n4586, Z => n1421);
   U5863 : AO2 port map( A => n4694, B => v_DATA_COLUMN_26_port, C => n4586, D 
                           => DATA_I(2), Z => n1422);
   U5864 : AO2 port map( A => n4694, B => v_DATA_COLUMN_25_port, C => DATA_I(1)
                           , D => n4586, Z => n1423);
   U5865 : AO2 port map( A => n4694, B => v_DATA_COLUMN_24_port, C => DATA_I(0)
                           , D => n4586, Z => n1424);
   U5866 : EON1 port map( A => n3956, B => n3704, C => VALID_DATA_I, D => n3704
                           , Z => n4312);
   U5867 : AO4 port map( A => CE_I, B => n4395, C => n4840, D => n1447, Z => 
                           n4346);
   U5868 : AO4 port map( A => n3948, B => n4713, C => n3947, D => CE_I, Z => 
                           n4301);
   U5869 : AO4 port map( A => n3949, B => n4713, C => n3948, D => CE_I, Z => 
                           n4302);
   U5870 : IVI port map( A => CE_I, Z => n4713);
   U5871 : IVI port map( A => RESET_I, Z => n4850);
   U5872 : IVI port map( A => n4356, Z => n4678);
   U5873 : IVI port map( A => n4355, Z => n4682);
   U5874 : IVI port map( A => n4357, Z => n4687);
   U5875 : IVI port map( A => n3359, Z => n4696);
   U5876 : IVI port map( A => n2957, Z => n4699);
   U5877 : IVI port map( A => n4361, Z => n4701);
   U5878 : IVI port map( A => n4359, Z => n4702);
   U5879 : IVI port map( A => n1959, Z => n4703);
   U5880 : IVI port map( A => n4379, Z => n4707);
   U5881 : IVI port map( A => n1609, Z => n4708);
   U5882 : IVI port map( A => n1527, Z => n4709);
   U5883 : IVI port map( A => n4349, Z => n4710);
   U5884 : IVA port map( A => n4496, Z => n4711);
   U5885 : ND2 port map( A => n4653, B => n4620, Z => n4714);
   U5886 : AO7 port map( A => n4620, B => n4653, C => n4714, Z => N199);
   U5887 : NR2 port map( A => n4714, B => v_INV_KEY_NUMB_2_port, Z => n4716);
   U5888 : AO6 port map( A => n4714, B => v_INV_KEY_NUMB_2_port, C => n4716, Z 
                           => n4715);
   U5889 : IV port map( A => n4715, Z => N200);
   U5890 : ND2 port map( A => n4716, B => n3942, Z => n4717);
   U5891 : AO7 port map( A => n4716, B => n3942, C => n4717, Z => N201);
   U5892 : EN port map( A => v_INV_KEY_NUMB_4_port, B => n4717, Z => N202);
   U5893 : NR2 port map( A => v_INV_KEY_NUMB_4_port, B => n4717, Z => n4718);
   U5894 : EO port map( A => v_INV_KEY_NUMB_5_port, B => n4718, Z => N203);
   U5895 : ND2 port map( A => v_CALCULATION_CNTR_1_port, B => 
                           v_CALCULATION_CNTR_0_port, Z => n4719);
   U5896 : EN port map( A => v_CALCULATION_CNTR_2_port, B => n4719, Z => N2084)
                           ;
   U5897 : AN3 port map( A => v_CALCULATION_CNTR_1_port, B => 
                           v_CALCULATION_CNTR_0_port, C => 
                           v_CALCULATION_CNTR_2_port, Z => n4721);
   U5898 : EO port map( A => v_CALCULATION_CNTR_3_port, B => n4721, Z => N2085)
                           ;
   U5899 : ND2 port map( A => v_CALCULATION_CNTR_3_port, B => n4721, Z => n4720
                           );
   U5900 : EN port map( A => v_CALCULATION_CNTR_4_port, B => n4720, Z => N2086)
                           ;
   U5901 : AN3 port map( A => v_CALCULATION_CNTR_3_port, B => n4721, C => 
                           v_CALCULATION_CNTR_4_port, Z => n4722);
   U5902 : EO port map( A => v_CALCULATION_CNTR_5_port, B => n4722, Z => N2087)
                           ;
   U5903 : ND2 port map( A => v_CALCULATION_CNTR_5_port, B => n4722, Z => n4723
                           );
   U5904 : EN port map( A => v_CALCULATION_CNTR_6_port, B => n4723, Z => N2088)
                           ;
   U5905 : NR2 port map( A => n4723, B => n4600, Z => n4724);
   U5906 : EO port map( A => v_CALCULATION_CNTR_7_port, B => n4724, Z => N2089)
                           ;
   U5907 : IVI port map( A => v_KEY_COLUMN_9_port, Z => n4725);
   U5908 : IVI port map( A => n449, Z => n4726);
   U5909 : IVI port map( A => n831, Z => n4727);
   U5910 : IVI port map( A => n459, Z => n4728);
   U5911 : IVI port map( A => n561, Z => n4729);
   U5912 : IVI port map( A => n551, Z => n4730);
   U5913 : IVI port map( A => n640, Z => n4731);
   U5914 : IVI port map( A => v_KEY_COLUMN_8_port, Z => n4732);
   U5915 : IVI port map( A => n995, Z => n4733);
   U5916 : IVI port map( A => n661, Z => n4734);
   U5917 : IVI port map( A => n766, Z => n4735);
   U5918 : IVI port map( A => n631, Z => n4736);
   U5919 : IVI port map( A => n781, Z => n4737);
   U5920 : IVI port map( A => n1289, Z => n4738);
   U5921 : IVI port map( A => n773, Z => n4739);
   U5922 : IVI port map( A => n639, Z => n4740);
   U5923 : IVI port map( A => n1364, Z => n4741);
   U5924 : IVI port map( A => n1102, Z => n4742);
   U5925 : IVI port map( A => n216, Z => n4743);
   U5926 : IVI port map( A => n224, Z => n4744);
   U5927 : IVI port map( A => n221, Z => n4745);
   U5928 : IVI port map( A => n1001, Z => n4746);
   U5929 : IVI port map( A => n1004, Z => n4747);
   U5930 : IVI port map( A => n1003, Z => n4748);
   U5931 : IVI port map( A => n1370, Z => n4749);
   U5932 : IVI port map( A => n1374, Z => n4750);
   U5933 : IVI port map( A => n1371, Z => n4751);
   U5934 : IVI port map( A => n231, Z => n4752);
   U5935 : IVI port map( A => n226, Z => n4753);
   U5936 : IVI port map( A => n202_port, Z => n4754);
   U5937 : IVI port map( A => n195, Z => n4755);
   U5938 : IVI port map( A => n1376, Z => n4756);
   U5939 : IVI port map( A => n423, Z => n4757);
   U5940 : IVI port map( A => n722, Z => n4758);
   U5941 : IVI port map( A => n729, Z => n4759);
   U5942 : IVI port map( A => v_KEY_COLUMN_4_port, Z => n4760);
   U5943 : IVI port map( A => v_KEY_COLUMN_3_port, Z => n4761);
   U5944 : IVI port map( A => n954, Z => n4762);
   U5945 : IVI port map( A => n964, Z => n4763);
   U5946 : IVI port map( A => n1100, Z => n4764);
   U5947 : IVI port map( A => n998, Z => n4765);
   U5948 : IVI port map( A => n673, Z => n4766);
   U5949 : IVI port map( A => n680, Z => n4767);
   U5950 : IVI port map( A => n1054, Z => n4768);
   U5951 : IVI port map( A => n1061, Z => n4769);
   U5952 : IVI port map( A => n192_port, Z => n4770);
   U5953 : IVI port map( A => v_KEY_COLUMN_2_port, Z => n4771);
   U5954 : IVI port map( A => n928, Z => n4772);
   U5955 : IVI port map( A => v_KEY_COLUMN_29_port, Z => n4773);
   U5956 : IVI port map( A => n1033, Z => n4774);
   U5957 : IVI port map( A => n850, Z => n4775);
   U5958 : IVI port map( A => n861, Z => n4776);
   U5959 : IVI port map( A => n866, Z => n4777);
   U5960 : IVI port map( A => n880, Z => n4778);
   U5961 : IVI port map( A => v_KEY_COLUMN_26_port, Z => n4779);
   U5962 : IVI port map( A => v_KEY_COLUMN_25_port, Z => n4780);
   U5963 : IVI port map( A => n827, Z => n4781);
   U5964 : IVI port map( A => n196, Z => n4782);
   U5965 : IVI port map( A => n182, Z => n4783);
   U5966 : IVI port map( A => n1997, Z => n4784);
   U5967 : IVI port map( A => v_KEY_COLUMN_21_port, Z => n4785);
   U5968 : IVI port map( A => n288, Z => n4786);
   U5969 : IVI port map( A => v_KEY_COLUMN_1_port, Z => n4787);
   U5970 : IVI port map( A => v_KEY_COLUMN_19_port, Z => n4788);
   U5971 : IVI port map( A => v_KEY_COLUMN_18_port, Z => n4789);
   U5972 : IVI port map( A => n121, Z => n4790);
   U5973 : IVI port map( A => n127, Z => n4791);
   U5974 : IVI port map( A => v_KEY_COLUMN_16_port, Z => n4792);
   U5975 : IVI port map( A => n179, Z => n4793);
   U5976 : IVI port map( A => n189, Z => n4794);
   U5977 : IVI port map( A => n402, Z => n4795);
   U5978 : IVI port map( A => n408, Z => n4796);
   U5979 : IVI port map( A => n414, Z => n4797);
   U5980 : IVI port map( A => n422, Z => n4798);
   U5981 : IVI port map( A => v_KEY_COLUMN_12_port, Z => n4799);
   U5982 : IVI port map( A => n338, Z => n4800);
   U5983 : IVI port map( A => n346, Z => n4801);
   U5984 : IVI port map( A => n352, Z => n4802);
   U5985 : IVI port map( A => n362, Z => n4803);
   U5986 : IVI port map( A => v_KEY_COLUMN_0_port, Z => n4804);
   U5987 : IVI port map( A => n157, Z => n4805);
   U5988 : IVI port map( A => n171, Z => n4806);
   U5989 : IVI port map( A => n656, Z => n4807);
   U5990 : IVI port map( A => n1407, Z => n4808);
   U5991 : IVI port map( A => n1414, Z => n4809);
   U5992 : IVI port map( A => n1426, Z => n4810);
   U5993 : IVI port map( A => n1437, Z => n4811);
   U5994 : IVI port map( A => n1410, Z => n4812);
   U5995 : IVI port map( A => n1417, Z => n4813);
   U5996 : IVI port map( A => n1429, Z => n4814);
   U5997 : IVI port map( A => n1438, Z => n4815);
   U5998 : IVI port map( A => n1411, Z => n4816);
   U5999 : IVI port map( A => n1419, Z => n4817);
   U6000 : IVI port map( A => n1430, Z => n4818);
   U6001 : IVI port map( A => n1439, Z => n4819);
   U6002 : IVI port map( A => n1412, Z => n4820);
   U6003 : IVI port map( A => n1420, Z => n4821);
   U6004 : IVI port map( A => n1431, Z => n4822);
   U6005 : IVI port map( A => n1440, Z => n4823);
   U6006 : IVI port map( A => n1413, Z => n4824);
   U6007 : IVI port map( A => n1421, Z => n4825);
   U6008 : IVI port map( A => n1433, Z => n4826);
   U6009 : IVI port map( A => n1441, Z => n4827);
   U6010 : IVI port map( A => n1418, Z => n4828);
   U6011 : IVI port map( A => n1422, Z => n4829);
   U6012 : IVI port map( A => n1434, Z => n4830);
   U6013 : IVI port map( A => n1442, Z => n4831);
   U6014 : IVI port map( A => n1403, Z => n4832);
   U6015 : IVI port map( A => n1423, Z => n4833);
   U6016 : IVI port map( A => n1432, Z => n4834);
   U6017 : IVI port map( A => n1435, Z => n4835);
   U6018 : IVI port map( A => n1406, Z => n4836);
   U6019 : IVI port map( A => n1424, Z => n4837);
   U6020 : IVI port map( A => n1436, Z => n4838);
   U6021 : IVI port map( A => n1443, Z => n4839);
   U6022 : IVI port map( A => VALID_DATA_I, Z => n4840);
   U6023 : IVI port map( A => n1398, Z => n4841);
   U6024 : IVI port map( A => n1486, Z => n4842);
   U6025 : IVI port map( A => n1487, Z => n4843);
   U6026 : IVI port map( A => n164, Z => n4844);
   U6027 : IVI port map( A => n1480, Z => n4845);
   U6028 : IVI port map( A => n1448, Z => n4846);
   U6029 : IVI port map( A => n1451, Z => n4847);
   U6030 : IVI port map( A => n1452, Z => n4848);
   U6031 : IVI port map( A => n1454, Z => n4849);
   U6032 : IVI port map( A => n1350, Z => n4851);
   U6033 : IVI port map( A => n1474, Z => n4852);
   U6034 : IVI port map( A => n1481, Z => n4853);
   U6035 : IVI port map( A => n1465, Z => n4854);
   U6036 : IVI port map( A => n103, Z => n4855);
   U6037 : IVI port map( A => n1353, Z => n4856);
   U6038 : IVI port map( A => n2391, Z => n4857);
   U6039 : IVI port map( A => n1509, Z => n4858);
   U6040 : IVI port map( A => n1485, Z => n4859);
   U6041 : IVI port map( A => n3672, Z => n4860);
   U6042 : IVI port map( A => n3802, Z => n4861);
   U6043 : IVI port map( A => n3798, Z => n4862);
   U6044 : IVI port map( A => n1498, Z => n4863);
   U6045 : IVI port map( A => n1499, Z => n4864);
   U6046 : IVI port map( A => n2813, Z => n4865);
   U6047 : IVI port map( A => n2606, Z => n4866);
   U6048 : IVI port map( A => n2792, Z => n4867);
   U6049 : IVI port map( A => n2560, Z => n4868);
   U6050 : IVI port map( A => n2677, Z => n4869);
   U6051 : IVI port map( A => n2639, Z => n4870);
   U6052 : IVI port map( A => n2713, Z => n4871);
   U6053 : IVI port map( A => n2850, Z => n4872);
   U6054 : IVI port map( A => n2635, Z => n4873);
   U6055 : IVI port map( A => n2871, Z => n4874);
   U6056 : IVI port map( A => n2692, Z => n4875);
   U6057 : IVI port map( A => n2719, Z => n4876);
   U6058 : IVI port map( A => n2653, Z => n4877);
   U6059 : IVI port map( A => n2542, Z => n4878);
   U6060 : IVI port map( A => n2874, Z => n4879);
   U6061 : IVI port map( A => n2591, Z => n4880);
   U6062 : IVI port map( A => n2738, Z => n4881);
   U6063 : IVI port map( A => n2528, Z => n4882);
   U6064 : IVI port map( A => n2529, Z => n4883);
   U6065 : IVI port map( A => n2540, Z => n4884);
   U6066 : IVI port map( A => n2649, Z => n4885);
   U6067 : IVI port map( A => n2678, Z => n4886);
   U6068 : IVI port map( A => n2803, Z => n4887);
   U6069 : IVI port map( A => n2728, Z => n4888);
   U6070 : IVI port map( A => n2532, Z => n4889);
   U6071 : IVI port map( A => n2587, Z => n4890);
   U6072 : IVI port map( A => n2583, Z => n4891);
   U6073 : IVI port map( A => n2562, Z => n4892);
   U6074 : IVI port map( A => n2624, Z => n4893);
   U6075 : IVI port map( A => n1955, Z => n4894);
   U6076 : IVI port map( A => n2715, Z => n4895);
   U6077 : IVI port map( A => n2714, Z => n4896);
   U6078 : IVI port map( A => n2507, Z => n4897);
   U6079 : IVI port map( A => n2676, Z => n4898);
   U6080 : IVI port map( A => n2739, Z => n4899);
   U6081 : IVI port map( A => n1988, Z => n4900);
   U6082 : IVI port map( A => n2549, Z => n4901);
   U6083 : IVI port map( A => n2568, Z => n4902);
   U6084 : IVI port map( A => n3043, Z => n4903);
   U6085 : IVI port map( A => n1868, Z => n4904);
   U6086 : IVI port map( A => n2333, Z => n4905);
   U6087 : IVI port map( A => n1897, Z => n4906);
   U6088 : IVI port map( A => n2294, Z => n4907);
   U6089 : IVI port map( A => n2413, Z => n4908);
   U6090 : IVI port map( A => n2074, Z => n4909);
   U6091 : IVI port map( A => n1912, Z => n4910);
   U6092 : IVI port map( A => n3445, Z => n4911);
   U6093 : IVI port map( A => n2665, Z => n4912);
   U6094 : IVI port map( A => n2590, Z => n4913);
   U6095 : IVI port map( A => n2584, Z => n4914);
   U6096 : IVI port map( A => n2550, Z => n4915);
   U6097 : IVI port map( A => n2759, Z => n4916);
   U6098 : IVI port map( A => n2965, Z => n4917);
   U6099 : IVI port map( A => n3053, Z => n4918);
   U6100 : IVI port map( A => n3057, Z => n4919);
   U6101 : IVI port map( A => n2963, Z => n4920);
   U6102 : IVI port map( A => n3083, Z => n4921);
   U6103 : IVI port map( A => n3210, Z => n4922);
   U6104 : IVI port map( A => n3288, Z => n4923);
   U6105 : IVI port map( A => n3285, Z => n4924);
   U6106 : IVI port map( A => n2987, Z => n4925);
   U6107 : IVI port map( A => n2953, Z => n4926);
   U6108 : IVI port map( A => n2970, Z => n4927);
   U6109 : IVI port map( A => n3221, Z => n4928);
   U6110 : IVI port map( A => n3132, Z => n4929);
   U6111 : IVI port map( A => n3200, Z => n4930);
   U6112 : IVI port map( A => n3097, Z => n4931);
   U6113 : IVI port map( A => n3123, Z => n4932);
   U6114 : IVI port map( A => n2993, Z => n4933);
   U6115 : IVI port map( A => n3118, Z => n4934);
   U6116 : IVI port map( A => n3070, Z => n4935);
   U6117 : IVI port map( A => n2990, Z => n4936);
   U6118 : IVI port map( A => n1688, Z => n4937);
   U6119 : IVI port map( A => n1722, Z => n4938);
   U6120 : IVI port map( A => n3119, Z => n4939);
   U6121 : IVI port map( A => n2947, Z => n4940);
   U6122 : IVI port map( A => n1713, Z => n4941);
   U6123 : IVI port map( A => n3142, Z => n4942);
   U6124 : IVI port map( A => n3143, Z => n4943);
   U6125 : IVI port map( A => n3254, Z => n4944);
   U6126 : IVI port map( A => n3009, Z => n4945);
   U6127 : IVI port map( A => n2954, Z => n4946);
   U6128 : IVI port map( A => n3117, Z => n4947);
   U6129 : IVI port map( A => n2986, Z => n4948);
   U6130 : IVI port map( A => n3182, Z => n4949);
   U6131 : IVI port map( A => n3039, Z => n4950);
   U6132 : IVI port map( A => n3007, Z => n4951);
   U6133 : IVI port map( A => n3163, Z => n4952);
   U6134 : IVI port map( A => n3081, Z => n4953);
   U6135 : IVI port map( A => n2933, Z => n4954);
   U6136 : IVI port map( A => n2094, Z => n4955);
   U6137 : IVI port map( A => n2190, Z => n4956);
   U6138 : IVI port map( A => n2341, Z => n4957);
   U6139 : IVI port map( A => n2372, Z => n4958);
   U6140 : IVI port map( A => n2158, Z => n4959);
   U6141 : IVI port map( A => n2072, Z => n4960);
   U6142 : IVI port map( A => n2133, Z => n4961);
   U6143 : IVI port map( A => n2087_port, Z => n4962);
   U6144 : IVI port map( A => n2347, Z => n4963);
   U6145 : IVI port map( A => n2064, Z => n4964);
   U6146 : IVI port map( A => n2130, Z => n4965);
   U6147 : IVI port map( A => n2154, Z => n4966);
   U6148 : IVI port map( A => n2066, Z => n4967);
   U6149 : IVI port map( A => n2236, Z => n4968);
   U6150 : IVI port map( A => n2159, Z => n4969);
   U6151 : IVI port map( A => n2178, Z => n4970);
   U6152 : IVI port map( A => n2153, Z => n4971);
   U6153 : IVI port map( A => n2162, Z => n4972);
   U6154 : IVI port map( A => n2239, Z => n4973);
   U6155 : IVI port map( A => n1916, Z => n4974);
   U6156 : IVI port map( A => n1900, Z => n4975);
   U6157 : IVI port map( A => n2044, Z => n4976);
   U6158 : IVI port map( A => n2306, Z => n4977);
   U6159 : IVI port map( A => n2120, Z => n4978);
   U6160 : IVI port map( A => n2038, Z => n4979);
   U6161 : IVI port map( A => n1914, Z => n4980);
   U6162 : IVI port map( A => n2095, Z => n4981);
   U6163 : IVI port map( A => n2380, Z => n4982);
   U6164 : IVI port map( A => n2075, Z => n4983);
   U6165 : IVI port map( A => n1906, Z => n4984);
   U6166 : IVI port map( A => n2261, Z => n4985);
   U6167 : IVI port map( A => n2084_port, Z => n4986);
   U6168 : IVI port map( A => n2121, Z => n4987);
   U6169 : IVI port map( A => n2165, Z => n4988);
   U6170 : IVI port map( A => n2344, Z => n4989);
   U6171 : IVI port map( A => n2186, Z => n4990);
   U6172 : IVI port map( A => n2245, Z => n4991);
   U6173 : IVI port map( A => n2128, Z => n4992);
   U6174 : IVI port map( A => n2060, Z => n4993);
   U6175 : IVI port map( A => n2408, Z => n4994);
   U6176 : IVI port map( A => n2047, Z => n4995);
   U6177 : IVI port map( A => n2129, Z => n4996);
   U6178 : IVI port map( A => n2281, Z => n4997);
   U6179 : IVI port map( A => n2227, Z => n4998);
   U6180 : IVI port map( A => n3367, Z => n4999);
   U6181 : IVI port map( A => n3455, Z => n5000);
   U6182 : IVI port map( A => n3459, Z => n5001);
   U6183 : IVI port map( A => n3365, Z => n5002);
   U6184 : IVI port map( A => n3485, Z => n5003);
   U6185 : IVI port map( A => n3611, Z => n5004);
   U6186 : IVI port map( A => n3692, Z => n5005);
   U6187 : IVI port map( A => n3689, Z => n5006);
   U6188 : IVI port map( A => n3388, Z => n5007);
   U6189 : IVI port map( A => n3355, Z => n5008);
   U6190 : IVI port map( A => n3372, Z => n5009);
   U6191 : IVI port map( A => n3622, Z => n5010);
   U6192 : IVI port map( A => n3533, Z => n5011);
   U6193 : IVI port map( A => n3601, Z => n5012);
   U6194 : IVI port map( A => n3499, Z => n5013);
   U6195 : IVI port map( A => n3524, Z => n5014);
   U6196 : IVI port map( A => n3394, Z => n5015);
   U6197 : IVI port map( A => n3519, Z => n5016);
   U6198 : IVI port map( A => n3472, Z => n5017);
   U6199 : IVI port map( A => n3391, Z => n5018);
   U6200 : IVI port map( A => n2454, Z => n5019);
   U6201 : IVI port map( A => n2486, Z => n5020);
   U6202 : IVI port map( A => n3520, Z => n5021);
   U6203 : IVI port map( A => n3349, Z => n5022);
   U6204 : IVI port map( A => n2477, Z => n5023);
   U6205 : IVI port map( A => n3543, Z => n5024);
   U6206 : IVI port map( A => n3544, Z => n5025);
   U6207 : IVI port map( A => n3656, Z => n5026);
   U6208 : IVI port map( A => n3410, Z => n5027);
   U6209 : IVI port map( A => n3356, Z => n5028);
   U6210 : IVI port map( A => n3518, Z => n5029);
   U6211 : IVI port map( A => n3387, Z => n5030);
   U6212 : IVI port map( A => n3583, Z => n5031);
   U6213 : IVI port map( A => n3440, Z => n5032);
   U6214 : IVI port map( A => n3408, Z => n5033);
   U6215 : IVI port map( A => n3564, Z => n5034);
   U6216 : IVI port map( A => n3483, Z => n5035);
   U6217 : IVI port map( A => n3335, Z => n5036);
   U6218 : IVI port map( A => n2946, Z => n5037);
   U6219 : IVI port map( A => n2949, Z => n5038);
   U6220 : IVI port map( A => n1877, Z => n5039);
   U6221 : IVI port map( A => n2541, Z => n5042);
   U6222 : IVI port map( A => n2544, Z => n5043);
   U6223 : IVI port map( A => n3348, Z => n5044);
   U6224 : IVI port map( A => n3351, Z => n5045);
   U6225 : IVI port map( A => n2476, Z => n5046);
   U6226 : IVI port map( A => n3342, Z => n5047);
   U6227 : IVI port map( A => n3325, Z => n5048);
   U6228 : IVI port map( A => n3338, Z => n5049);
   U6229 : IVI port map( A => n3389, Z => n5050);
   U6230 : IVI port map( A => n3457, Z => n5051);
   U6231 : IVI port map( A => n1712, Z => n5052);
   U6232 : IVI port map( A => n2940, Z => n5053);
   U6233 : IVI port map( A => n2923, Z => n5054);
   U6234 : IVI port map( A => n2936, Z => n5055);
   U6235 : IVI port map( A => n2988, Z => n5056);
   U6236 : IVI port map( A => n3055, Z => n5057);
   U6237 : IVI port map( A => n1978, Z => n5058);
   U6238 : IVI port map( A => n2585, Z => n5059);
   U6239 : IVI port map( A => n2651, Z => n5060);
   U6240 : IVI port map( A => n2534, Z => n5061);
   U6241 : IVI port map( A => n2519, Z => n5062);
   U6242 : IVI port map( A => n2530, Z => n5063);
   U6243 : IVI port map( A => n1901, Z => n5064);
   U6244 : IVI port map( A => n2935, Z => n5065);
   U6245 : IVI port map( A => n2911, Z => n5066);
   U6246 : IVI port map( A => n3082, Z => n5067);
   U6247 : IVI port map( A => n3027, Z => n5068);
   U6248 : IVI port map( A => n2093, Z => n5069);
   U6249 : IVI port map( A => n3337, Z => n5070);
   U6250 : IVI port map( A => n3313, Z => n5071);
   U6251 : IVI port map( A => n3484, Z => n5072);
   U6252 : IVI port map( A => n3428, Z => n5073);

end SYN_Behavioral;
